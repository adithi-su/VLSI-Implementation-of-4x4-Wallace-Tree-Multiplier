magic
tech scmos
timestamp 1636353112
<< nwell >>
rect 0 1276 17 1325
rect 139 1246 171 1263
rect 0 1189 17 1238
rect 77 1223 109 1240
rect 197 1236 229 1253
rect 367 1247 399 1264
rect 305 1224 337 1241
rect 425 1237 457 1254
rect 139 1197 171 1214
rect 207 1192 227 1208
rect 367 1198 399 1215
rect 435 1193 455 1209
rect 1 1101 18 1150
rect 2 1020 19 1069
rect 126 992 158 1009
rect 2 936 19 985
rect 64 969 96 986
rect 184 982 216 999
rect 306 992 338 1009
rect 244 969 276 986
rect 364 982 396 999
rect 621 989 653 1006
rect 559 966 591 983
rect 679 979 711 996
rect 126 943 158 960
rect 194 938 214 954
rect 306 943 338 960
rect 374 938 394 954
rect 407 946 456 961
rect 621 940 653 957
rect 689 935 709 951
rect 2 849 19 898
rect 329 821 361 838
rect 3 761 20 810
rect 267 798 299 815
rect 387 811 419 828
rect 509 821 541 838
rect 447 798 479 815
rect 567 811 599 828
rect 329 772 361 789
rect 397 767 417 783
rect 509 772 541 789
rect 577 767 597 783
rect 609 775 658 790
rect 4 680 21 729
rect 124 654 156 671
rect 4 596 21 645
rect 62 631 94 648
rect 182 644 214 661
rect 304 654 336 671
rect 242 631 274 648
rect 362 644 394 661
rect 657 656 689 673
rect 595 633 627 650
rect 715 646 747 663
rect 837 656 869 673
rect 775 633 807 650
rect 895 646 927 663
rect 124 605 156 622
rect 192 600 212 616
rect 304 605 336 622
rect 372 600 392 616
rect 405 608 454 623
rect 657 607 689 624
rect 725 602 745 618
rect 837 607 869 624
rect 905 602 925 618
rect 937 610 986 625
rect 4 509 21 558
rect 315 499 347 516
rect 253 476 285 493
rect 373 489 405 506
rect 495 499 527 516
rect 433 476 465 493
rect 553 489 585 506
rect 5 421 22 470
rect 315 450 347 467
rect 383 445 403 461
rect 495 450 527 467
rect 563 445 583 461
rect 595 453 644 468
rect 145 398 177 415
rect 6 340 23 389
rect 83 375 115 392
rect 203 388 235 405
rect 145 349 177 366
rect 562 364 594 381
rect 213 344 233 360
rect 500 341 532 358
rect 620 354 652 371
rect 742 364 774 381
rect 680 341 712 358
rect 800 354 832 371
rect 562 315 594 332
rect 630 310 650 326
rect 742 315 774 332
rect 810 310 830 326
rect 842 318 891 333
rect 6 256 23 305
rect 6 169 23 218
rect 162 212 194 229
rect 100 189 132 206
rect 220 202 252 219
rect 342 212 374 229
rect 280 189 312 206
rect 400 202 432 219
rect 162 163 194 180
rect 230 158 250 174
rect 342 163 374 180
rect 410 158 430 174
rect 442 166 491 181
rect 585 165 617 182
rect 523 142 555 159
rect 643 155 675 172
rect 765 165 797 182
rect 703 142 735 159
rect 823 155 855 172
rect 7 81 24 130
rect 585 116 617 133
rect 653 111 673 127
rect 765 116 797 133
rect 833 111 853 127
rect 865 119 914 134
rect 8 0 25 49
<< polysilicon >>
rect 7 1317 9 1319
rect 15 1318 32 1319
rect 15 1317 17 1318
rect 21 1317 32 1318
rect 35 1317 38 1319
rect 7 1301 9 1303
rect 15 1302 32 1303
rect 15 1301 24 1302
rect 28 1301 32 1302
rect 35 1301 37 1303
rect 7 1281 9 1283
rect 15 1282 32 1283
rect 15 1281 17 1282
rect 21 1281 32 1282
rect 35 1281 37 1283
rect 144 1254 146 1256
rect 164 1254 166 1256
rect 372 1255 374 1257
rect 392 1255 394 1257
rect 144 1246 146 1248
rect 145 1242 146 1246
rect 7 1230 9 1232
rect 15 1231 32 1232
rect 15 1230 17 1231
rect 21 1230 32 1231
rect 35 1230 38 1232
rect 82 1231 84 1233
rect 102 1231 104 1233
rect 144 1231 146 1242
rect 164 1239 166 1248
rect 372 1247 374 1249
rect 202 1244 204 1246
rect 222 1244 224 1246
rect 165 1235 166 1239
rect 373 1243 374 1247
rect 202 1236 204 1238
rect 164 1231 166 1235
rect 203 1232 204 1236
rect 144 1226 146 1228
rect 164 1226 166 1228
rect 82 1223 84 1225
rect 83 1219 84 1223
rect 7 1214 9 1216
rect 15 1215 32 1216
rect 15 1214 24 1215
rect 28 1214 32 1215
rect 35 1214 37 1216
rect 82 1208 84 1219
rect 102 1216 104 1225
rect 202 1221 204 1232
rect 222 1229 224 1238
rect 310 1232 312 1234
rect 330 1232 332 1234
rect 223 1225 224 1229
rect 372 1232 374 1243
rect 392 1240 394 1249
rect 430 1245 432 1247
rect 450 1245 452 1247
rect 393 1236 394 1240
rect 430 1237 432 1239
rect 392 1232 394 1236
rect 431 1233 432 1237
rect 372 1227 374 1229
rect 392 1227 394 1229
rect 222 1221 224 1225
rect 310 1224 312 1226
rect 311 1220 312 1224
rect 202 1216 204 1218
rect 222 1216 224 1218
rect 103 1212 104 1216
rect 102 1208 104 1212
rect 144 1205 146 1207
rect 164 1205 166 1207
rect 82 1203 84 1205
rect 102 1203 104 1205
rect 310 1209 312 1220
rect 330 1217 332 1226
rect 430 1222 432 1233
rect 450 1230 452 1239
rect 451 1226 452 1230
rect 450 1222 452 1226
rect 430 1217 432 1219
rect 450 1217 452 1219
rect 331 1213 332 1217
rect 330 1209 332 1213
rect 372 1206 374 1208
rect 392 1206 394 1208
rect 310 1204 312 1206
rect 330 1204 332 1206
rect 215 1199 217 1201
rect 443 1200 445 1202
rect 144 1197 146 1199
rect 7 1194 9 1196
rect 15 1195 32 1196
rect 15 1194 17 1195
rect 21 1194 32 1195
rect 35 1194 37 1196
rect 145 1193 146 1197
rect 144 1182 146 1193
rect 164 1190 166 1199
rect 372 1198 374 1200
rect 373 1194 374 1198
rect 215 1190 217 1193
rect 165 1186 166 1190
rect 164 1182 166 1186
rect 215 1182 217 1186
rect 144 1177 146 1179
rect 164 1177 166 1179
rect 215 1177 217 1179
rect 372 1183 374 1194
rect 392 1191 394 1200
rect 443 1191 445 1194
rect 393 1187 394 1191
rect 392 1183 394 1187
rect 443 1183 445 1187
rect 372 1178 374 1180
rect 392 1178 394 1180
rect 443 1178 445 1180
rect 8 1142 10 1144
rect 16 1143 33 1144
rect 16 1142 18 1143
rect 22 1142 33 1143
rect 36 1142 39 1144
rect 8 1126 10 1128
rect 16 1127 33 1128
rect 16 1126 25 1127
rect 29 1126 33 1127
rect 36 1126 38 1128
rect 8 1106 10 1108
rect 16 1107 33 1108
rect 16 1106 18 1107
rect 22 1106 33 1107
rect 36 1106 38 1108
rect 9 1061 11 1063
rect 17 1062 34 1063
rect 17 1061 19 1062
rect 23 1061 34 1062
rect 37 1061 40 1063
rect 9 1045 11 1047
rect 17 1046 34 1047
rect 17 1045 26 1046
rect 30 1045 34 1046
rect 37 1045 39 1047
rect 9 1025 11 1027
rect 17 1026 34 1027
rect 17 1025 19 1026
rect 23 1025 34 1026
rect 37 1025 39 1027
rect 131 1000 133 1002
rect 151 1000 153 1002
rect 311 1000 313 1002
rect 331 1000 333 1002
rect 626 997 628 999
rect 646 997 648 999
rect 131 992 133 994
rect 132 988 133 992
rect 9 977 11 979
rect 17 978 34 979
rect 17 977 19 978
rect 23 977 34 978
rect 37 977 40 979
rect 69 977 71 979
rect 89 977 91 979
rect 131 977 133 988
rect 151 985 153 994
rect 311 992 313 994
rect 189 990 191 992
rect 209 990 211 992
rect 152 981 153 985
rect 312 988 313 992
rect 189 982 191 984
rect 151 977 153 981
rect 190 978 191 982
rect 131 972 133 974
rect 151 972 153 974
rect 69 969 71 971
rect 70 965 71 969
rect 9 961 11 963
rect 17 962 34 963
rect 17 961 26 962
rect 30 961 34 962
rect 37 961 39 963
rect 69 954 71 965
rect 89 962 91 971
rect 189 967 191 978
rect 209 975 211 984
rect 249 977 251 979
rect 269 977 271 979
rect 210 971 211 975
rect 311 977 313 988
rect 331 985 333 994
rect 369 990 371 992
rect 389 990 391 992
rect 332 981 333 985
rect 626 989 628 991
rect 627 985 628 989
rect 369 982 371 984
rect 331 977 333 981
rect 370 978 371 982
rect 311 972 313 974
rect 331 972 333 974
rect 209 967 211 971
rect 249 969 251 971
rect 250 965 251 969
rect 189 962 191 964
rect 209 962 211 964
rect 90 958 91 962
rect 89 954 91 958
rect 131 951 133 953
rect 151 951 153 953
rect 69 949 71 951
rect 89 949 91 951
rect 249 954 251 965
rect 269 962 271 971
rect 369 967 371 978
rect 389 975 391 984
rect 390 971 391 975
rect 564 974 566 976
rect 584 974 586 976
rect 389 967 391 971
rect 626 974 628 985
rect 646 982 648 991
rect 684 987 686 989
rect 704 987 706 989
rect 647 978 648 982
rect 684 979 686 981
rect 646 974 648 978
rect 685 975 686 979
rect 626 969 628 971
rect 646 969 648 971
rect 564 966 566 968
rect 369 962 371 964
rect 389 962 391 964
rect 565 962 566 966
rect 270 958 271 962
rect 269 954 271 958
rect 311 951 313 953
rect 331 951 333 953
rect 249 949 251 951
rect 269 949 271 951
rect 202 945 204 947
rect 412 953 414 955
rect 428 953 430 955
rect 448 953 450 955
rect 564 951 566 962
rect 584 959 586 968
rect 684 964 686 975
rect 704 972 706 981
rect 705 968 706 972
rect 704 964 706 968
rect 684 959 686 961
rect 704 959 706 961
rect 585 955 586 959
rect 584 951 586 955
rect 626 948 628 950
rect 646 948 648 950
rect 382 945 384 947
rect 131 943 133 945
rect 9 941 11 943
rect 17 942 34 943
rect 17 941 19 942
rect 23 941 34 942
rect 37 941 39 943
rect 132 939 133 943
rect 131 928 133 939
rect 151 936 153 945
rect 311 943 313 945
rect 312 939 313 943
rect 202 936 204 939
rect 152 932 153 936
rect 151 928 153 932
rect 202 928 204 932
rect 131 923 133 925
rect 151 923 153 925
rect 202 923 204 925
rect 311 928 313 939
rect 331 936 333 945
rect 382 936 384 939
rect 332 932 333 936
rect 412 935 414 947
rect 428 944 430 947
rect 429 940 430 944
rect 331 928 333 932
rect 382 928 384 932
rect 413 931 414 935
rect 311 923 313 925
rect 331 923 333 925
rect 382 923 384 925
rect 412 927 414 931
rect 428 927 430 940
rect 448 935 450 947
rect 564 946 566 948
rect 584 946 586 948
rect 697 942 699 944
rect 626 940 628 942
rect 627 936 628 940
rect 448 928 450 931
rect 412 922 414 924
rect 428 922 430 924
rect 448 922 450 924
rect 626 925 628 936
rect 646 933 648 942
rect 697 933 699 936
rect 647 929 648 933
rect 646 925 648 929
rect 697 925 699 929
rect 626 920 628 922
rect 646 920 648 922
rect 697 920 699 922
rect 9 890 11 892
rect 17 891 34 892
rect 17 890 19 891
rect 23 890 34 891
rect 37 890 40 892
rect 9 874 11 876
rect 17 875 34 876
rect 17 874 26 875
rect 30 874 34 875
rect 37 874 39 876
rect 9 854 11 856
rect 17 855 34 856
rect 17 854 19 855
rect 23 854 34 855
rect 37 854 39 856
rect 334 829 336 831
rect 354 829 356 831
rect 514 829 516 831
rect 534 829 536 831
rect 334 821 336 823
rect 335 817 336 821
rect 272 806 274 808
rect 292 806 294 808
rect 10 802 12 804
rect 18 803 35 804
rect 18 802 20 803
rect 24 802 35 803
rect 38 802 41 804
rect 334 806 336 817
rect 354 814 356 823
rect 514 821 516 823
rect 392 819 394 821
rect 412 819 414 821
rect 355 810 356 814
rect 515 817 516 821
rect 392 811 394 813
rect 354 806 356 810
rect 393 807 394 811
rect 334 801 336 803
rect 354 801 356 803
rect 272 798 274 800
rect 273 794 274 798
rect 10 786 12 788
rect 18 787 35 788
rect 18 786 27 787
rect 31 786 35 787
rect 38 786 40 788
rect 272 783 274 794
rect 292 791 294 800
rect 392 796 394 807
rect 412 804 414 813
rect 452 806 454 808
rect 472 806 474 808
rect 413 800 414 804
rect 514 806 516 817
rect 534 814 536 823
rect 572 819 574 821
rect 592 819 594 821
rect 535 810 536 814
rect 572 811 574 813
rect 534 806 536 810
rect 573 807 574 811
rect 514 801 516 803
rect 534 801 536 803
rect 412 796 414 800
rect 452 798 454 800
rect 453 794 454 798
rect 392 791 394 793
rect 412 791 414 793
rect 293 787 294 791
rect 292 783 294 787
rect 334 780 336 782
rect 354 780 356 782
rect 272 778 274 780
rect 292 778 294 780
rect 452 783 454 794
rect 472 791 474 800
rect 572 796 574 807
rect 592 804 594 813
rect 593 800 594 804
rect 592 796 594 800
rect 572 791 574 793
rect 592 791 594 793
rect 473 787 474 791
rect 472 783 474 787
rect 514 780 516 782
rect 534 780 536 782
rect 452 778 454 780
rect 472 778 474 780
rect 405 774 407 776
rect 614 782 616 784
rect 630 782 632 784
rect 650 782 652 784
rect 585 774 587 776
rect 334 772 336 774
rect 335 768 336 772
rect 10 766 12 768
rect 18 767 35 768
rect 18 766 20 767
rect 24 766 35 767
rect 38 766 40 768
rect 334 757 336 768
rect 354 765 356 774
rect 514 772 516 774
rect 515 768 516 772
rect 405 765 407 768
rect 355 761 356 765
rect 354 757 356 761
rect 405 757 407 761
rect 334 752 336 754
rect 354 752 356 754
rect 405 752 407 754
rect 514 757 516 768
rect 534 765 536 774
rect 585 765 587 768
rect 535 761 536 765
rect 614 764 616 776
rect 630 773 632 776
rect 631 769 632 773
rect 534 757 536 761
rect 585 757 587 761
rect 615 760 616 764
rect 514 752 516 754
rect 534 752 536 754
rect 585 752 587 754
rect 614 756 616 760
rect 630 756 632 769
rect 650 764 652 776
rect 650 757 652 760
rect 614 751 616 753
rect 630 751 632 753
rect 650 751 652 753
rect 11 721 13 723
rect 19 722 36 723
rect 19 721 21 722
rect 25 721 36 722
rect 39 721 42 723
rect 11 705 13 707
rect 19 706 36 707
rect 19 705 28 706
rect 32 705 36 706
rect 39 705 41 707
rect 11 685 13 687
rect 19 686 36 687
rect 19 685 21 686
rect 25 685 36 686
rect 39 685 41 687
rect 662 664 664 666
rect 682 664 684 666
rect 842 664 844 666
rect 862 664 864 666
rect 129 662 131 664
rect 149 662 151 664
rect 309 662 311 664
rect 329 662 331 664
rect 662 656 664 658
rect 129 654 131 656
rect 130 650 131 654
rect 67 639 69 641
rect 87 639 89 641
rect 11 637 13 639
rect 19 638 36 639
rect 19 637 21 638
rect 25 637 36 638
rect 39 637 42 639
rect 129 639 131 650
rect 149 647 151 656
rect 309 654 311 656
rect 187 652 189 654
rect 207 652 209 654
rect 150 643 151 647
rect 310 650 311 654
rect 187 644 189 646
rect 149 639 151 643
rect 188 640 189 644
rect 129 634 131 636
rect 149 634 151 636
rect 67 631 69 633
rect 68 627 69 631
rect 11 621 13 623
rect 19 622 36 623
rect 19 621 28 622
rect 32 621 36 622
rect 39 621 41 623
rect 67 616 69 627
rect 87 624 89 633
rect 187 629 189 640
rect 207 637 209 646
rect 247 639 249 641
rect 267 639 269 641
rect 208 633 209 637
rect 309 639 311 650
rect 329 647 331 656
rect 367 652 369 654
rect 387 652 389 654
rect 663 652 664 656
rect 330 643 331 647
rect 367 644 369 646
rect 329 639 331 643
rect 368 640 369 644
rect 309 634 311 636
rect 329 634 331 636
rect 207 629 209 633
rect 247 631 249 633
rect 248 627 249 631
rect 187 624 189 626
rect 207 624 209 626
rect 88 620 89 624
rect 87 616 89 620
rect 129 613 131 615
rect 149 613 151 615
rect 67 611 69 613
rect 87 611 89 613
rect 247 616 249 627
rect 267 624 269 633
rect 367 629 369 640
rect 387 637 389 646
rect 600 641 602 643
rect 620 641 622 643
rect 388 633 389 637
rect 662 641 664 652
rect 682 649 684 658
rect 842 656 844 658
rect 720 654 722 656
rect 740 654 742 656
rect 683 645 684 649
rect 843 652 844 656
rect 720 646 722 648
rect 682 641 684 645
rect 721 642 722 646
rect 662 636 664 638
rect 682 636 684 638
rect 600 633 602 635
rect 387 629 389 633
rect 601 629 602 633
rect 367 624 369 626
rect 387 624 389 626
rect 268 620 269 624
rect 267 616 269 620
rect 309 613 311 615
rect 329 613 331 615
rect 247 611 249 613
rect 267 611 269 613
rect 200 607 202 609
rect 410 615 412 617
rect 426 615 428 617
rect 446 615 448 617
rect 600 618 602 629
rect 620 626 622 635
rect 720 631 722 642
rect 740 639 742 648
rect 780 641 782 643
rect 800 641 802 643
rect 741 635 742 639
rect 842 641 844 652
rect 862 649 864 658
rect 900 654 902 656
rect 920 654 922 656
rect 863 645 864 649
rect 900 646 902 648
rect 862 641 864 645
rect 901 642 902 646
rect 842 636 844 638
rect 862 636 864 638
rect 740 631 742 635
rect 780 633 782 635
rect 781 629 782 633
rect 720 626 722 628
rect 740 626 742 628
rect 621 622 622 626
rect 620 618 622 622
rect 662 615 664 617
rect 682 615 684 617
rect 600 613 602 615
rect 620 613 622 615
rect 780 618 782 629
rect 800 626 802 635
rect 900 631 902 642
rect 920 639 922 648
rect 921 635 922 639
rect 920 631 922 635
rect 900 626 902 628
rect 920 626 922 628
rect 801 622 802 626
rect 800 618 802 622
rect 842 615 844 617
rect 862 615 864 617
rect 780 613 782 615
rect 800 613 802 615
rect 733 609 735 611
rect 942 617 944 619
rect 958 617 960 619
rect 978 617 980 619
rect 913 609 915 611
rect 380 607 382 609
rect 129 605 131 607
rect 11 601 13 603
rect 19 602 36 603
rect 19 601 21 602
rect 25 601 36 602
rect 39 601 41 603
rect 130 601 131 605
rect 129 590 131 601
rect 149 598 151 607
rect 309 605 311 607
rect 310 601 311 605
rect 200 598 202 601
rect 150 594 151 598
rect 149 590 151 594
rect 200 590 202 594
rect 129 585 131 587
rect 149 585 151 587
rect 200 585 202 587
rect 309 590 311 601
rect 329 598 331 607
rect 380 598 382 601
rect 330 594 331 598
rect 410 597 412 609
rect 426 606 428 609
rect 427 602 428 606
rect 329 590 331 594
rect 380 590 382 594
rect 411 593 412 597
rect 309 585 311 587
rect 329 585 331 587
rect 380 585 382 587
rect 410 589 412 593
rect 426 589 428 602
rect 446 597 448 609
rect 662 607 664 609
rect 663 603 664 607
rect 446 590 448 593
rect 662 592 664 603
rect 682 600 684 609
rect 842 607 844 609
rect 843 603 844 607
rect 733 600 735 603
rect 683 596 684 600
rect 682 592 684 596
rect 733 592 735 596
rect 662 587 664 589
rect 682 587 684 589
rect 733 587 735 589
rect 842 592 844 603
rect 862 600 864 609
rect 913 600 915 603
rect 863 596 864 600
rect 942 599 944 611
rect 958 608 960 611
rect 959 604 960 608
rect 862 592 864 596
rect 913 592 915 596
rect 943 595 944 599
rect 842 587 844 589
rect 862 587 864 589
rect 913 587 915 589
rect 942 591 944 595
rect 958 591 960 604
rect 978 599 980 611
rect 978 592 980 595
rect 942 586 944 588
rect 958 586 960 588
rect 978 586 980 588
rect 410 584 412 586
rect 426 584 428 586
rect 446 584 448 586
rect 11 550 13 552
rect 19 551 36 552
rect 19 550 21 551
rect 25 550 36 551
rect 39 550 42 552
rect 11 534 13 536
rect 19 535 36 536
rect 19 534 28 535
rect 32 534 36 535
rect 39 534 41 536
rect 11 514 13 516
rect 19 515 36 516
rect 19 514 21 515
rect 25 514 36 515
rect 39 514 41 516
rect 320 507 322 509
rect 340 507 342 509
rect 500 507 502 509
rect 520 507 522 509
rect 320 499 322 501
rect 321 495 322 499
rect 258 484 260 486
rect 278 484 280 486
rect 320 484 322 495
rect 340 492 342 501
rect 500 499 502 501
rect 378 497 380 499
rect 398 497 400 499
rect 341 488 342 492
rect 501 495 502 499
rect 378 489 380 491
rect 340 484 342 488
rect 379 485 380 489
rect 320 479 322 481
rect 340 479 342 481
rect 258 476 260 478
rect 259 472 260 476
rect 12 462 14 464
rect 20 463 37 464
rect 20 462 22 463
rect 26 462 37 463
rect 40 462 43 464
rect 258 461 260 472
rect 278 469 280 478
rect 378 474 380 485
rect 398 482 400 491
rect 438 484 440 486
rect 458 484 460 486
rect 399 478 400 482
rect 500 484 502 495
rect 520 492 522 501
rect 558 497 560 499
rect 578 497 580 499
rect 521 488 522 492
rect 558 489 560 491
rect 520 484 522 488
rect 559 485 560 489
rect 500 479 502 481
rect 520 479 522 481
rect 398 474 400 478
rect 438 476 440 478
rect 439 472 440 476
rect 378 469 380 471
rect 398 469 400 471
rect 279 465 280 469
rect 278 461 280 465
rect 320 458 322 460
rect 340 458 342 460
rect 258 456 260 458
rect 278 456 280 458
rect 438 461 440 472
rect 458 469 460 478
rect 558 474 560 485
rect 578 482 580 491
rect 579 478 580 482
rect 578 474 580 478
rect 558 469 560 471
rect 578 469 580 471
rect 459 465 460 469
rect 458 461 460 465
rect 500 458 502 460
rect 520 458 522 460
rect 438 456 440 458
rect 458 456 460 458
rect 391 452 393 454
rect 600 460 602 462
rect 616 460 618 462
rect 636 460 638 462
rect 571 452 573 454
rect 320 450 322 452
rect 12 446 14 448
rect 20 447 37 448
rect 20 446 29 447
rect 33 446 37 447
rect 40 446 42 448
rect 321 446 322 450
rect 320 435 322 446
rect 340 443 342 452
rect 500 450 502 452
rect 501 446 502 450
rect 391 443 393 446
rect 341 439 342 443
rect 340 435 342 439
rect 391 435 393 439
rect 320 430 322 432
rect 340 430 342 432
rect 391 430 393 432
rect 500 435 502 446
rect 520 443 522 452
rect 571 443 573 446
rect 521 439 522 443
rect 600 442 602 454
rect 616 451 618 454
rect 617 447 618 451
rect 520 435 522 439
rect 571 435 573 439
rect 601 438 602 442
rect 500 430 502 432
rect 520 430 522 432
rect 571 430 573 432
rect 600 434 602 438
rect 616 434 618 447
rect 636 442 638 454
rect 636 435 638 438
rect 600 429 602 431
rect 616 429 618 431
rect 636 429 638 431
rect 12 426 14 428
rect 20 427 37 428
rect 20 426 22 427
rect 26 426 37 427
rect 40 426 42 428
rect 150 406 152 408
rect 170 406 172 408
rect 150 398 152 400
rect 151 394 152 398
rect 88 383 90 385
rect 108 383 110 385
rect 13 381 15 383
rect 21 382 38 383
rect 21 381 23 382
rect 27 381 38 382
rect 41 381 44 383
rect 150 383 152 394
rect 170 391 172 400
rect 208 396 210 398
rect 228 396 230 398
rect 171 387 172 391
rect 208 388 210 390
rect 170 383 172 387
rect 209 384 210 388
rect 150 378 152 380
rect 170 378 172 380
rect 88 375 90 377
rect 89 371 90 375
rect 13 365 15 367
rect 21 366 38 367
rect 21 365 30 366
rect 34 365 38 366
rect 41 365 43 367
rect 88 360 90 371
rect 108 368 110 377
rect 208 373 210 384
rect 228 381 230 390
rect 229 377 230 381
rect 228 373 230 377
rect 567 372 569 374
rect 587 372 589 374
rect 747 372 749 374
rect 767 372 769 374
rect 208 368 210 370
rect 228 368 230 370
rect 109 364 110 368
rect 108 360 110 364
rect 567 364 569 366
rect 568 360 569 364
rect 150 357 152 359
rect 170 357 172 359
rect 88 355 90 357
rect 108 355 110 357
rect 221 351 223 353
rect 150 349 152 351
rect 13 345 15 347
rect 21 346 38 347
rect 21 345 23 346
rect 27 345 38 346
rect 41 345 43 347
rect 151 345 152 349
rect 150 334 152 345
rect 170 342 172 351
rect 505 349 507 351
rect 525 349 527 351
rect 221 342 223 345
rect 567 349 569 360
rect 587 357 589 366
rect 747 364 749 366
rect 625 362 627 364
rect 645 362 647 364
rect 588 353 589 357
rect 748 360 749 364
rect 625 354 627 356
rect 587 349 589 353
rect 626 350 627 354
rect 567 344 569 346
rect 587 344 589 346
rect 171 338 172 342
rect 505 341 507 343
rect 170 334 172 338
rect 221 334 223 338
rect 506 337 507 341
rect 150 329 152 331
rect 170 329 172 331
rect 221 329 223 331
rect 505 326 507 337
rect 525 334 527 343
rect 625 339 627 350
rect 645 347 647 356
rect 685 349 687 351
rect 705 349 707 351
rect 646 343 647 347
rect 747 349 749 360
rect 767 357 769 366
rect 805 362 807 364
rect 825 362 827 364
rect 768 353 769 357
rect 805 354 807 356
rect 767 349 769 353
rect 806 350 807 354
rect 747 344 749 346
rect 767 344 769 346
rect 645 339 647 343
rect 685 341 687 343
rect 686 337 687 341
rect 625 334 627 336
rect 645 334 647 336
rect 526 330 527 334
rect 525 326 527 330
rect 567 323 569 325
rect 587 323 589 325
rect 505 321 507 323
rect 525 321 527 323
rect 685 326 687 337
rect 705 334 707 343
rect 805 339 807 350
rect 825 347 827 356
rect 826 343 827 347
rect 825 339 827 343
rect 805 334 807 336
rect 825 334 827 336
rect 706 330 707 334
rect 705 326 707 330
rect 747 323 749 325
rect 767 323 769 325
rect 685 321 687 323
rect 705 321 707 323
rect 638 317 640 319
rect 847 325 849 327
rect 863 325 865 327
rect 883 325 885 327
rect 818 317 820 319
rect 567 315 569 317
rect 568 311 569 315
rect 13 297 15 299
rect 21 298 38 299
rect 21 297 23 298
rect 27 297 38 298
rect 41 297 44 299
rect 567 300 569 311
rect 587 308 589 317
rect 747 315 749 317
rect 748 311 749 315
rect 638 308 640 311
rect 588 304 589 308
rect 587 300 589 304
rect 638 300 640 304
rect 567 295 569 297
rect 587 295 589 297
rect 638 295 640 297
rect 747 300 749 311
rect 767 308 769 317
rect 818 308 820 311
rect 768 304 769 308
rect 847 307 849 319
rect 863 316 865 319
rect 864 312 865 316
rect 767 300 769 304
rect 818 300 820 304
rect 848 303 849 307
rect 747 295 749 297
rect 767 295 769 297
rect 818 295 820 297
rect 847 299 849 303
rect 863 299 865 312
rect 883 307 885 319
rect 883 300 885 303
rect 847 294 849 296
rect 863 294 865 296
rect 883 294 885 296
rect 13 281 15 283
rect 21 282 38 283
rect 21 281 30 282
rect 34 281 38 282
rect 41 281 43 283
rect 13 261 15 263
rect 21 262 38 263
rect 21 261 23 262
rect 27 261 38 262
rect 41 261 43 263
rect 167 220 169 222
rect 187 220 189 222
rect 347 220 349 222
rect 367 220 369 222
rect 167 212 169 214
rect 13 210 15 212
rect 21 211 38 212
rect 21 210 23 211
rect 27 210 38 211
rect 41 210 44 212
rect 168 208 169 212
rect 105 197 107 199
rect 125 197 127 199
rect 13 194 15 196
rect 21 195 38 196
rect 21 194 30 195
rect 34 194 38 195
rect 41 194 43 196
rect 167 197 169 208
rect 187 205 189 214
rect 347 212 349 214
rect 225 210 227 212
rect 245 210 247 212
rect 188 201 189 205
rect 348 208 349 212
rect 225 202 227 204
rect 187 197 189 201
rect 226 198 227 202
rect 167 192 169 194
rect 187 192 189 194
rect 105 189 107 191
rect 106 185 107 189
rect 13 174 15 176
rect 21 175 38 176
rect 21 174 23 175
rect 27 174 38 175
rect 41 174 43 176
rect 105 174 107 185
rect 125 182 127 191
rect 225 187 227 198
rect 245 195 247 204
rect 285 197 287 199
rect 305 197 307 199
rect 246 191 247 195
rect 347 197 349 208
rect 367 205 369 214
rect 405 210 407 212
rect 425 210 427 212
rect 368 201 369 205
rect 405 202 407 204
rect 367 197 369 201
rect 406 198 407 202
rect 347 192 349 194
rect 367 192 369 194
rect 245 187 247 191
rect 285 189 287 191
rect 286 185 287 189
rect 225 182 227 184
rect 245 182 247 184
rect 126 178 127 182
rect 125 174 127 178
rect 167 171 169 173
rect 187 171 189 173
rect 105 169 107 171
rect 125 169 127 171
rect 285 174 287 185
rect 305 182 307 191
rect 405 187 407 198
rect 425 195 427 204
rect 426 191 427 195
rect 425 187 427 191
rect 405 182 407 184
rect 425 182 427 184
rect 306 178 307 182
rect 305 174 307 178
rect 347 171 349 173
rect 367 171 369 173
rect 285 169 287 171
rect 305 169 307 171
rect 238 165 240 167
rect 447 173 449 175
rect 463 173 465 175
rect 483 173 485 175
rect 590 173 592 175
rect 610 173 612 175
rect 770 173 772 175
rect 790 173 792 175
rect 418 165 420 167
rect 167 163 169 165
rect 168 159 169 163
rect 167 148 169 159
rect 187 156 189 165
rect 347 163 349 165
rect 348 159 349 163
rect 238 156 240 159
rect 188 152 189 156
rect 187 148 189 152
rect 238 148 240 152
rect 167 143 169 145
rect 187 143 189 145
rect 238 143 240 145
rect 347 148 349 159
rect 367 156 369 165
rect 418 156 420 159
rect 368 152 369 156
rect 447 155 449 167
rect 463 164 465 167
rect 464 160 465 164
rect 367 148 369 152
rect 418 148 420 152
rect 448 151 449 155
rect 347 143 349 145
rect 367 143 369 145
rect 418 143 420 145
rect 447 147 449 151
rect 463 147 465 160
rect 483 155 485 167
rect 590 165 592 167
rect 591 161 592 165
rect 483 148 485 151
rect 528 150 530 152
rect 548 150 550 152
rect 590 150 592 161
rect 610 158 612 167
rect 770 165 772 167
rect 648 163 650 165
rect 668 163 670 165
rect 611 154 612 158
rect 771 161 772 165
rect 648 155 650 157
rect 610 150 612 154
rect 649 151 650 155
rect 590 145 592 147
rect 610 145 612 147
rect 447 142 449 144
rect 463 142 465 144
rect 483 142 485 144
rect 528 142 530 144
rect 529 138 530 142
rect 528 127 530 138
rect 548 135 550 144
rect 648 140 650 151
rect 668 148 670 157
rect 708 150 710 152
rect 728 150 730 152
rect 669 144 670 148
rect 770 150 772 161
rect 790 158 792 167
rect 828 163 830 165
rect 848 163 850 165
rect 791 154 792 158
rect 828 155 830 157
rect 790 150 792 154
rect 829 151 830 155
rect 770 145 772 147
rect 790 145 792 147
rect 668 140 670 144
rect 708 142 710 144
rect 709 138 710 142
rect 648 135 650 137
rect 668 135 670 137
rect 549 131 550 135
rect 548 127 550 131
rect 590 124 592 126
rect 610 124 612 126
rect 14 122 16 124
rect 22 123 39 124
rect 22 122 24 123
rect 28 122 39 123
rect 42 122 45 124
rect 528 122 530 124
rect 548 122 550 124
rect 708 127 710 138
rect 728 135 730 144
rect 828 140 830 151
rect 848 148 850 157
rect 849 144 850 148
rect 848 140 850 144
rect 828 135 830 137
rect 848 135 850 137
rect 729 131 730 135
rect 728 127 730 131
rect 770 124 772 126
rect 790 124 792 126
rect 708 122 710 124
rect 728 122 730 124
rect 661 118 663 120
rect 870 126 872 128
rect 886 126 888 128
rect 906 126 908 128
rect 841 118 843 120
rect 590 116 592 118
rect 591 112 592 116
rect 14 106 16 108
rect 22 107 39 108
rect 22 106 31 107
rect 35 106 39 107
rect 42 106 44 108
rect 590 101 592 112
rect 610 109 612 118
rect 770 116 772 118
rect 771 112 772 116
rect 661 109 663 112
rect 611 105 612 109
rect 610 101 612 105
rect 661 101 663 105
rect 590 96 592 98
rect 610 96 612 98
rect 661 96 663 98
rect 770 101 772 112
rect 790 109 792 118
rect 841 109 843 112
rect 791 105 792 109
rect 870 108 872 120
rect 886 117 888 120
rect 887 113 888 117
rect 790 101 792 105
rect 841 101 843 105
rect 871 104 872 108
rect 770 96 772 98
rect 790 96 792 98
rect 841 96 843 98
rect 870 100 872 104
rect 886 100 888 113
rect 906 108 908 120
rect 906 101 908 104
rect 870 95 872 97
rect 886 95 888 97
rect 906 95 908 97
rect 14 86 16 88
rect 22 87 39 88
rect 22 86 24 87
rect 28 86 39 87
rect 42 86 44 88
rect 15 41 17 43
rect 23 42 40 43
rect 23 41 25 42
rect 29 41 40 42
rect 43 41 46 43
rect 15 25 17 27
rect 23 26 40 27
rect 23 25 32 26
rect 36 25 40 26
rect 43 25 45 27
rect 15 5 17 7
rect 23 6 40 7
rect 23 5 25 6
rect 29 5 40 6
rect 43 5 45 7
<< ndiffusion >>
rect 32 1319 35 1320
rect 32 1316 35 1317
rect 32 1303 35 1304
rect 32 1283 35 1301
rect 32 1280 35 1281
rect 32 1232 35 1233
rect 32 1229 35 1230
rect 143 1228 144 1231
rect 146 1228 164 1231
rect 166 1228 167 1231
rect 32 1216 35 1217
rect 32 1196 35 1214
rect 371 1229 372 1232
rect 374 1229 392 1232
rect 394 1229 395 1232
rect 201 1218 202 1221
rect 204 1218 222 1221
rect 224 1218 225 1221
rect 81 1205 82 1208
rect 84 1205 102 1208
rect 104 1205 105 1208
rect 429 1219 430 1222
rect 432 1219 450 1222
rect 452 1219 453 1222
rect 309 1206 310 1209
rect 312 1206 330 1209
rect 332 1206 333 1209
rect 32 1193 35 1194
rect 143 1179 144 1182
rect 146 1179 164 1182
rect 166 1179 167 1182
rect 213 1179 215 1182
rect 217 1179 219 1182
rect 371 1180 372 1183
rect 374 1180 392 1183
rect 394 1180 395 1183
rect 441 1180 443 1183
rect 445 1180 447 1183
rect 33 1144 36 1145
rect 33 1141 36 1142
rect 33 1128 36 1129
rect 33 1108 36 1126
rect 33 1105 36 1106
rect 34 1063 37 1064
rect 34 1060 37 1061
rect 34 1047 37 1048
rect 34 1027 37 1045
rect 34 1024 37 1025
rect 34 979 37 980
rect 34 976 37 977
rect 130 974 131 977
rect 133 974 151 977
rect 153 974 154 977
rect 34 963 37 964
rect 34 943 37 961
rect 310 974 311 977
rect 313 974 331 977
rect 333 974 334 977
rect 188 964 189 967
rect 191 964 209 967
rect 211 964 212 967
rect 68 951 69 954
rect 71 951 89 954
rect 91 951 92 954
rect 625 971 626 974
rect 628 971 646 974
rect 648 971 649 974
rect 368 964 369 967
rect 371 964 389 967
rect 391 964 392 967
rect 248 951 249 954
rect 251 951 269 954
rect 271 951 272 954
rect 683 961 684 964
rect 686 961 704 964
rect 706 961 707 964
rect 563 948 564 951
rect 566 948 584 951
rect 586 948 587 951
rect 34 940 37 941
rect 130 925 131 928
rect 133 925 151 928
rect 153 925 154 928
rect 200 925 202 928
rect 204 925 206 928
rect 310 925 311 928
rect 313 925 331 928
rect 333 925 334 928
rect 380 925 382 928
rect 384 925 386 928
rect 411 924 412 927
rect 414 924 415 927
rect 427 924 428 927
rect 430 924 431 927
rect 446 924 448 928
rect 450 924 452 928
rect 625 922 626 925
rect 628 922 646 925
rect 648 922 649 925
rect 695 922 697 925
rect 699 922 701 925
rect 34 892 37 893
rect 34 889 37 890
rect 34 876 37 877
rect 34 856 37 874
rect 34 853 37 854
rect 35 804 38 805
rect 35 801 38 802
rect 333 803 334 806
rect 336 803 354 806
rect 356 803 357 806
rect 35 788 38 789
rect 35 768 38 786
rect 513 803 514 806
rect 516 803 534 806
rect 536 803 537 806
rect 391 793 392 796
rect 394 793 412 796
rect 414 793 415 796
rect 271 780 272 783
rect 274 780 292 783
rect 294 780 295 783
rect 571 793 572 796
rect 574 793 592 796
rect 594 793 595 796
rect 451 780 452 783
rect 454 780 472 783
rect 474 780 475 783
rect 35 765 38 766
rect 333 754 334 757
rect 336 754 354 757
rect 356 754 357 757
rect 403 754 405 757
rect 407 754 409 757
rect 513 754 514 757
rect 516 754 534 757
rect 536 754 537 757
rect 583 754 585 757
rect 587 754 589 757
rect 613 753 614 756
rect 616 753 617 756
rect 629 753 630 756
rect 632 753 633 756
rect 648 753 650 757
rect 652 753 654 757
rect 36 723 39 724
rect 36 720 39 721
rect 36 707 39 708
rect 36 687 39 705
rect 36 684 39 685
rect 36 639 39 640
rect 36 636 39 637
rect 128 636 129 639
rect 131 636 149 639
rect 151 636 152 639
rect 36 623 39 624
rect 36 603 39 621
rect 308 636 309 639
rect 311 636 329 639
rect 331 636 332 639
rect 186 626 187 629
rect 189 626 207 629
rect 209 626 210 629
rect 66 613 67 616
rect 69 613 87 616
rect 89 613 90 616
rect 661 638 662 641
rect 664 638 682 641
rect 684 638 685 641
rect 366 626 367 629
rect 369 626 387 629
rect 389 626 390 629
rect 246 613 247 616
rect 249 613 267 616
rect 269 613 270 616
rect 841 638 842 641
rect 844 638 862 641
rect 864 638 865 641
rect 719 628 720 631
rect 722 628 740 631
rect 742 628 743 631
rect 599 615 600 618
rect 602 615 620 618
rect 622 615 623 618
rect 899 628 900 631
rect 902 628 920 631
rect 922 628 923 631
rect 779 615 780 618
rect 782 615 800 618
rect 802 615 803 618
rect 36 600 39 601
rect 128 587 129 590
rect 131 587 149 590
rect 151 587 152 590
rect 198 587 200 590
rect 202 587 204 590
rect 308 587 309 590
rect 311 587 329 590
rect 331 587 332 590
rect 378 587 380 590
rect 382 587 384 590
rect 409 586 410 589
rect 412 586 413 589
rect 425 586 426 589
rect 428 586 429 589
rect 444 586 446 590
rect 448 586 450 590
rect 661 589 662 592
rect 664 589 682 592
rect 684 589 685 592
rect 731 589 733 592
rect 735 589 737 592
rect 841 589 842 592
rect 844 589 862 592
rect 864 589 865 592
rect 911 589 913 592
rect 915 589 917 592
rect 941 588 942 591
rect 944 588 945 591
rect 957 588 958 591
rect 960 588 961 591
rect 976 588 978 592
rect 980 588 982 592
rect 36 552 39 553
rect 36 549 39 550
rect 36 536 39 537
rect 36 516 39 534
rect 36 513 39 514
rect 319 481 320 484
rect 322 481 340 484
rect 342 481 343 484
rect 37 464 40 465
rect 37 461 40 462
rect 499 481 500 484
rect 502 481 520 484
rect 522 481 523 484
rect 377 471 378 474
rect 380 471 398 474
rect 400 471 401 474
rect 257 458 258 461
rect 260 458 278 461
rect 280 458 281 461
rect 557 471 558 474
rect 560 471 578 474
rect 580 471 581 474
rect 437 458 438 461
rect 440 458 458 461
rect 460 458 461 461
rect 37 448 40 449
rect 37 428 40 446
rect 319 432 320 435
rect 322 432 340 435
rect 342 432 343 435
rect 389 432 391 435
rect 393 432 395 435
rect 499 432 500 435
rect 502 432 520 435
rect 522 432 523 435
rect 569 432 571 435
rect 573 432 575 435
rect 599 431 600 434
rect 602 431 603 434
rect 615 431 616 434
rect 618 431 619 434
rect 634 431 636 435
rect 638 431 640 435
rect 37 425 40 426
rect 38 383 41 384
rect 38 380 41 381
rect 149 380 150 383
rect 152 380 170 383
rect 172 380 173 383
rect 38 367 41 368
rect 38 347 41 365
rect 207 370 208 373
rect 210 370 228 373
rect 230 370 231 373
rect 87 357 88 360
rect 90 357 108 360
rect 110 357 111 360
rect 38 344 41 345
rect 566 346 567 349
rect 569 346 587 349
rect 589 346 590 349
rect 149 331 150 334
rect 152 331 170 334
rect 172 331 173 334
rect 219 331 221 334
rect 223 331 225 334
rect 746 346 747 349
rect 749 346 767 349
rect 769 346 770 349
rect 624 336 625 339
rect 627 336 645 339
rect 647 336 648 339
rect 504 323 505 326
rect 507 323 525 326
rect 527 323 528 326
rect 804 336 805 339
rect 807 336 825 339
rect 827 336 828 339
rect 684 323 685 326
rect 687 323 705 326
rect 707 323 708 326
rect 38 299 41 300
rect 566 297 567 300
rect 569 297 587 300
rect 589 297 590 300
rect 38 296 41 297
rect 636 297 638 300
rect 640 297 642 300
rect 746 297 747 300
rect 749 297 767 300
rect 769 297 770 300
rect 816 297 818 300
rect 820 297 822 300
rect 846 296 847 299
rect 849 296 850 299
rect 862 296 863 299
rect 865 296 866 299
rect 881 296 883 300
rect 885 296 887 300
rect 38 283 41 284
rect 38 263 41 281
rect 38 260 41 261
rect 38 212 41 213
rect 38 209 41 210
rect 38 196 41 197
rect 38 176 41 194
rect 166 194 167 197
rect 169 194 187 197
rect 189 194 190 197
rect 38 173 41 174
rect 346 194 347 197
rect 349 194 367 197
rect 369 194 370 197
rect 224 184 225 187
rect 227 184 245 187
rect 247 184 248 187
rect 104 171 105 174
rect 107 171 125 174
rect 127 171 128 174
rect 404 184 405 187
rect 407 184 425 187
rect 427 184 428 187
rect 284 171 285 174
rect 287 171 305 174
rect 307 171 308 174
rect 166 145 167 148
rect 169 145 187 148
rect 189 145 190 148
rect 236 145 238 148
rect 240 145 242 148
rect 346 145 347 148
rect 349 145 367 148
rect 369 145 370 148
rect 416 145 418 148
rect 420 145 422 148
rect 446 144 447 147
rect 449 144 450 147
rect 462 144 463 147
rect 465 144 466 147
rect 481 144 483 148
rect 485 144 487 148
rect 589 147 590 150
rect 592 147 610 150
rect 612 147 613 150
rect 39 124 42 125
rect 769 147 770 150
rect 772 147 790 150
rect 792 147 793 150
rect 647 137 648 140
rect 650 137 668 140
rect 670 137 671 140
rect 527 124 528 127
rect 530 124 548 127
rect 550 124 551 127
rect 39 121 42 122
rect 827 137 828 140
rect 830 137 848 140
rect 850 137 851 140
rect 707 124 708 127
rect 710 124 728 127
rect 730 124 731 127
rect 39 108 42 109
rect 39 88 42 106
rect 589 98 590 101
rect 592 98 610 101
rect 612 98 613 101
rect 659 98 661 101
rect 663 98 665 101
rect 769 98 770 101
rect 772 98 790 101
rect 792 98 793 101
rect 839 98 841 101
rect 843 98 845 101
rect 869 97 870 100
rect 872 97 873 100
rect 885 97 886 100
rect 888 97 889 100
rect 904 97 906 101
rect 908 97 910 101
rect 39 85 42 86
rect 40 43 43 44
rect 40 40 43 41
rect 40 27 43 28
rect 40 7 43 25
rect 40 4 43 5
<< pdiffusion >>
rect 9 1321 10 1323
rect 14 1321 15 1323
rect 9 1319 15 1321
rect 9 1316 15 1317
rect 9 1313 10 1316
rect 14 1313 15 1316
rect 9 1304 10 1306
rect 14 1304 15 1306
rect 9 1303 15 1304
rect 9 1300 15 1301
rect 9 1298 10 1300
rect 14 1298 15 1300
rect 9 1284 10 1286
rect 14 1284 15 1286
rect 9 1283 15 1284
rect 9 1280 15 1281
rect 9 1278 10 1280
rect 14 1278 15 1280
rect 369 1254 372 1255
rect 141 1253 144 1254
rect 143 1249 144 1253
rect 141 1248 144 1249
rect 146 1253 149 1254
rect 161 1253 164 1254
rect 146 1249 147 1253
rect 163 1249 164 1253
rect 146 1248 149 1249
rect 161 1248 164 1249
rect 166 1253 169 1254
rect 166 1249 167 1253
rect 371 1250 372 1254
rect 369 1249 372 1250
rect 374 1254 377 1255
rect 389 1254 392 1255
rect 374 1250 375 1254
rect 391 1250 392 1254
rect 374 1249 377 1250
rect 389 1249 392 1250
rect 394 1254 397 1255
rect 394 1250 395 1254
rect 394 1249 397 1250
rect 166 1248 169 1249
rect 9 1234 10 1236
rect 14 1234 15 1236
rect 9 1232 15 1234
rect 9 1229 15 1230
rect 9 1226 10 1229
rect 14 1226 15 1229
rect 79 1230 82 1231
rect 81 1226 82 1230
rect 79 1225 82 1226
rect 84 1230 87 1231
rect 99 1230 102 1231
rect 84 1226 85 1230
rect 101 1226 102 1230
rect 84 1225 87 1226
rect 99 1225 102 1226
rect 104 1230 107 1231
rect 104 1226 105 1230
rect 199 1243 202 1244
rect 201 1239 202 1243
rect 199 1238 202 1239
rect 204 1243 207 1244
rect 219 1243 222 1244
rect 204 1239 205 1243
rect 221 1239 222 1243
rect 204 1238 207 1239
rect 219 1238 222 1239
rect 224 1243 227 1244
rect 224 1239 225 1243
rect 224 1238 227 1239
rect 104 1225 107 1226
rect 9 1217 10 1219
rect 14 1217 15 1219
rect 9 1216 15 1217
rect 9 1213 15 1214
rect 9 1211 10 1213
rect 14 1211 15 1213
rect 9 1197 10 1199
rect 14 1197 15 1199
rect 9 1196 15 1197
rect 307 1231 310 1232
rect 309 1227 310 1231
rect 307 1226 310 1227
rect 312 1231 315 1232
rect 327 1231 330 1232
rect 312 1227 313 1231
rect 329 1227 330 1231
rect 312 1226 315 1227
rect 327 1226 330 1227
rect 332 1231 335 1232
rect 332 1227 333 1231
rect 427 1244 430 1245
rect 429 1240 430 1244
rect 427 1239 430 1240
rect 432 1244 435 1245
rect 447 1244 450 1245
rect 432 1240 433 1244
rect 449 1240 450 1244
rect 432 1239 435 1240
rect 447 1239 450 1240
rect 452 1244 455 1245
rect 452 1240 453 1244
rect 452 1239 455 1240
rect 332 1226 335 1227
rect 141 1204 144 1205
rect 143 1200 144 1204
rect 141 1199 144 1200
rect 146 1204 149 1205
rect 161 1204 164 1205
rect 146 1200 147 1204
rect 163 1200 164 1204
rect 146 1199 149 1200
rect 161 1199 164 1200
rect 166 1204 169 1205
rect 369 1205 372 1206
rect 166 1200 167 1204
rect 371 1201 372 1205
rect 166 1199 169 1200
rect 369 1200 372 1201
rect 374 1205 377 1206
rect 389 1205 392 1206
rect 374 1201 375 1205
rect 391 1201 392 1205
rect 374 1200 377 1201
rect 389 1200 392 1201
rect 394 1205 397 1206
rect 394 1201 395 1205
rect 394 1200 397 1201
rect 9 1193 15 1194
rect 9 1191 10 1193
rect 14 1191 15 1193
rect 212 1198 215 1199
rect 214 1194 215 1198
rect 212 1193 215 1194
rect 217 1198 221 1199
rect 217 1194 218 1198
rect 217 1193 221 1194
rect 440 1199 443 1200
rect 442 1195 443 1199
rect 440 1194 443 1195
rect 445 1199 449 1200
rect 445 1195 446 1199
rect 445 1194 449 1195
rect 10 1146 11 1148
rect 15 1146 16 1148
rect 10 1144 16 1146
rect 10 1141 16 1142
rect 10 1138 11 1141
rect 15 1138 16 1141
rect 10 1129 11 1131
rect 15 1129 16 1131
rect 10 1128 16 1129
rect 10 1125 16 1126
rect 10 1123 11 1125
rect 15 1123 16 1125
rect 10 1109 11 1111
rect 15 1109 16 1111
rect 10 1108 16 1109
rect 10 1105 16 1106
rect 10 1103 11 1105
rect 15 1103 16 1105
rect 11 1065 12 1067
rect 16 1065 17 1067
rect 11 1063 17 1065
rect 11 1060 17 1061
rect 11 1057 12 1060
rect 16 1057 17 1060
rect 11 1048 12 1050
rect 16 1048 17 1050
rect 11 1047 17 1048
rect 11 1044 17 1045
rect 11 1042 12 1044
rect 16 1042 17 1044
rect 11 1028 12 1030
rect 16 1028 17 1030
rect 11 1027 17 1028
rect 11 1024 17 1025
rect 11 1022 12 1024
rect 16 1022 17 1024
rect 128 999 131 1000
rect 130 995 131 999
rect 128 994 131 995
rect 133 999 136 1000
rect 148 999 151 1000
rect 133 995 134 999
rect 150 995 151 999
rect 133 994 136 995
rect 148 994 151 995
rect 153 999 156 1000
rect 308 999 311 1000
rect 153 995 154 999
rect 310 995 311 999
rect 153 994 156 995
rect 308 994 311 995
rect 313 999 316 1000
rect 328 999 331 1000
rect 313 995 314 999
rect 330 995 331 999
rect 313 994 316 995
rect 328 994 331 995
rect 333 999 336 1000
rect 333 995 334 999
rect 623 996 626 997
rect 333 994 336 995
rect 11 981 12 983
rect 16 981 17 983
rect 11 979 17 981
rect 11 976 17 977
rect 11 973 12 976
rect 16 973 17 976
rect 66 976 69 977
rect 68 972 69 976
rect 66 971 69 972
rect 71 976 74 977
rect 86 976 89 977
rect 71 972 72 976
rect 88 972 89 976
rect 71 971 74 972
rect 86 971 89 972
rect 91 976 94 977
rect 91 972 92 976
rect 186 989 189 990
rect 188 985 189 989
rect 186 984 189 985
rect 191 989 194 990
rect 206 989 209 990
rect 191 985 192 989
rect 208 985 209 989
rect 191 984 194 985
rect 206 984 209 985
rect 211 989 214 990
rect 211 985 212 989
rect 211 984 214 985
rect 91 971 94 972
rect 11 964 12 966
rect 16 964 17 966
rect 11 963 17 964
rect 11 960 17 961
rect 11 958 12 960
rect 16 958 17 960
rect 11 944 12 946
rect 16 944 17 946
rect 11 943 17 944
rect 246 976 249 977
rect 248 972 249 976
rect 246 971 249 972
rect 251 976 254 977
rect 266 976 269 977
rect 251 972 252 976
rect 268 972 269 976
rect 251 971 254 972
rect 266 971 269 972
rect 271 976 274 977
rect 271 972 272 976
rect 625 992 626 996
rect 623 991 626 992
rect 628 996 631 997
rect 643 996 646 997
rect 628 992 629 996
rect 645 992 646 996
rect 628 991 631 992
rect 643 991 646 992
rect 648 996 651 997
rect 648 992 649 996
rect 648 991 651 992
rect 366 989 369 990
rect 368 985 369 989
rect 366 984 369 985
rect 371 989 374 990
rect 386 989 389 990
rect 371 985 372 989
rect 388 985 389 989
rect 371 984 374 985
rect 386 984 389 985
rect 391 989 394 990
rect 391 985 392 989
rect 391 984 394 985
rect 271 971 274 972
rect 128 950 131 951
rect 130 946 131 950
rect 128 945 131 946
rect 133 950 136 951
rect 148 950 151 951
rect 133 946 134 950
rect 150 946 151 950
rect 133 945 136 946
rect 148 945 151 946
rect 153 950 156 951
rect 561 973 564 974
rect 563 969 564 973
rect 561 968 564 969
rect 566 973 569 974
rect 581 973 584 974
rect 566 969 567 973
rect 583 969 584 973
rect 566 968 569 969
rect 581 968 584 969
rect 586 973 589 974
rect 586 969 587 973
rect 681 986 684 987
rect 683 982 684 986
rect 681 981 684 982
rect 686 986 689 987
rect 701 986 704 987
rect 686 982 687 986
rect 703 982 704 986
rect 686 981 689 982
rect 701 981 704 982
rect 706 986 709 987
rect 706 982 707 986
rect 706 981 709 982
rect 586 968 589 969
rect 153 946 154 950
rect 308 950 311 951
rect 153 945 156 946
rect 310 946 311 950
rect 308 945 311 946
rect 313 950 316 951
rect 328 950 331 951
rect 313 946 314 950
rect 330 946 331 950
rect 313 945 316 946
rect 328 945 331 946
rect 333 950 336 951
rect 409 952 412 953
rect 333 946 334 950
rect 411 948 412 952
rect 409 947 412 948
rect 414 947 428 953
rect 430 952 434 953
rect 443 952 448 953
rect 430 948 431 952
rect 446 948 448 952
rect 430 947 434 948
rect 443 947 448 948
rect 450 952 455 953
rect 450 948 452 952
rect 450 947 455 948
rect 333 945 336 946
rect 11 940 17 941
rect 11 938 12 940
rect 16 938 17 940
rect 199 944 202 945
rect 201 940 202 944
rect 199 939 202 940
rect 204 944 208 945
rect 204 940 205 944
rect 204 939 208 940
rect 379 944 382 945
rect 381 940 382 944
rect 379 939 382 940
rect 384 944 388 945
rect 384 940 385 944
rect 384 939 388 940
rect 623 947 626 948
rect 625 943 626 947
rect 623 942 626 943
rect 628 947 631 948
rect 643 947 646 948
rect 628 943 629 947
rect 645 943 646 947
rect 628 942 631 943
rect 643 942 646 943
rect 648 947 651 948
rect 648 943 649 947
rect 648 942 651 943
rect 694 941 697 942
rect 696 937 697 941
rect 694 936 697 937
rect 699 941 703 942
rect 699 937 700 941
rect 699 936 703 937
rect 11 894 12 896
rect 16 894 17 896
rect 11 892 17 894
rect 11 889 17 890
rect 11 886 12 889
rect 16 886 17 889
rect 11 877 12 879
rect 16 877 17 879
rect 11 876 17 877
rect 11 873 17 874
rect 11 871 12 873
rect 16 871 17 873
rect 11 857 12 859
rect 16 857 17 859
rect 11 856 17 857
rect 11 853 17 854
rect 11 851 12 853
rect 16 851 17 853
rect 331 828 334 829
rect 333 824 334 828
rect 331 823 334 824
rect 336 828 339 829
rect 351 828 354 829
rect 336 824 337 828
rect 353 824 354 828
rect 336 823 339 824
rect 351 823 354 824
rect 356 828 359 829
rect 511 828 514 829
rect 356 824 357 828
rect 513 824 514 828
rect 356 823 359 824
rect 511 823 514 824
rect 516 828 519 829
rect 531 828 534 829
rect 516 824 517 828
rect 533 824 534 828
rect 516 823 519 824
rect 531 823 534 824
rect 536 828 539 829
rect 536 824 537 828
rect 536 823 539 824
rect 12 806 13 808
rect 17 806 18 808
rect 12 804 18 806
rect 269 805 272 806
rect 12 801 18 802
rect 12 798 13 801
rect 17 798 18 801
rect 271 801 272 805
rect 269 800 272 801
rect 274 805 277 806
rect 289 805 292 806
rect 274 801 275 805
rect 291 801 292 805
rect 274 800 277 801
rect 289 800 292 801
rect 294 805 297 806
rect 294 801 295 805
rect 389 818 392 819
rect 391 814 392 818
rect 389 813 392 814
rect 394 818 397 819
rect 409 818 412 819
rect 394 814 395 818
rect 411 814 412 818
rect 394 813 397 814
rect 409 813 412 814
rect 414 818 417 819
rect 414 814 415 818
rect 414 813 417 814
rect 294 800 297 801
rect 12 789 13 791
rect 17 789 18 791
rect 12 788 18 789
rect 12 785 18 786
rect 12 783 13 785
rect 17 783 18 785
rect 12 769 13 771
rect 17 769 18 771
rect 12 768 18 769
rect 449 805 452 806
rect 451 801 452 805
rect 449 800 452 801
rect 454 805 457 806
rect 469 805 472 806
rect 454 801 455 805
rect 471 801 472 805
rect 454 800 457 801
rect 469 800 472 801
rect 474 805 477 806
rect 474 801 475 805
rect 569 818 572 819
rect 571 814 572 818
rect 569 813 572 814
rect 574 818 577 819
rect 589 818 592 819
rect 574 814 575 818
rect 591 814 592 818
rect 574 813 577 814
rect 589 813 592 814
rect 594 818 597 819
rect 594 814 595 818
rect 594 813 597 814
rect 474 800 477 801
rect 331 779 334 780
rect 333 775 334 779
rect 331 774 334 775
rect 336 779 339 780
rect 351 779 354 780
rect 336 775 337 779
rect 353 775 354 779
rect 336 774 339 775
rect 351 774 354 775
rect 356 779 359 780
rect 356 775 357 779
rect 511 779 514 780
rect 356 774 359 775
rect 513 775 514 779
rect 511 774 514 775
rect 516 779 519 780
rect 531 779 534 780
rect 516 775 517 779
rect 533 775 534 779
rect 516 774 519 775
rect 531 774 534 775
rect 536 779 539 780
rect 611 781 614 782
rect 536 775 537 779
rect 613 777 614 781
rect 611 776 614 777
rect 616 776 630 782
rect 632 781 636 782
rect 645 781 650 782
rect 632 777 633 781
rect 648 777 650 781
rect 632 776 636 777
rect 645 776 650 777
rect 652 781 657 782
rect 652 777 654 781
rect 652 776 657 777
rect 536 774 539 775
rect 12 765 18 766
rect 12 763 13 765
rect 17 763 18 765
rect 402 773 405 774
rect 404 769 405 773
rect 402 768 405 769
rect 407 773 411 774
rect 407 769 408 773
rect 407 768 411 769
rect 582 773 585 774
rect 584 769 585 773
rect 582 768 585 769
rect 587 773 591 774
rect 587 769 588 773
rect 587 768 591 769
rect 13 725 14 727
rect 18 725 19 727
rect 13 723 19 725
rect 13 720 19 721
rect 13 717 14 720
rect 18 717 19 720
rect 13 708 14 710
rect 18 708 19 710
rect 13 707 19 708
rect 13 704 19 705
rect 13 702 14 704
rect 18 702 19 704
rect 13 688 14 690
rect 18 688 19 690
rect 13 687 19 688
rect 13 684 19 685
rect 13 682 14 684
rect 18 682 19 684
rect 659 663 662 664
rect 126 661 129 662
rect 128 657 129 661
rect 126 656 129 657
rect 131 661 134 662
rect 146 661 149 662
rect 131 657 132 661
rect 148 657 149 661
rect 131 656 134 657
rect 146 656 149 657
rect 151 661 154 662
rect 306 661 309 662
rect 151 657 152 661
rect 308 657 309 661
rect 151 656 154 657
rect 306 656 309 657
rect 311 661 314 662
rect 326 661 329 662
rect 311 657 312 661
rect 328 657 329 661
rect 311 656 314 657
rect 326 656 329 657
rect 331 661 334 662
rect 331 657 332 661
rect 661 659 662 663
rect 659 658 662 659
rect 664 663 667 664
rect 679 663 682 664
rect 664 659 665 663
rect 681 659 682 663
rect 664 658 667 659
rect 679 658 682 659
rect 684 663 687 664
rect 839 663 842 664
rect 684 659 685 663
rect 841 659 842 663
rect 684 658 687 659
rect 839 658 842 659
rect 844 663 847 664
rect 859 663 862 664
rect 844 659 845 663
rect 861 659 862 663
rect 844 658 847 659
rect 859 658 862 659
rect 864 663 867 664
rect 864 659 865 663
rect 864 658 867 659
rect 331 656 334 657
rect 13 641 14 643
rect 18 641 19 643
rect 13 639 19 641
rect 13 636 19 637
rect 13 633 14 636
rect 18 633 19 636
rect 64 638 67 639
rect 66 634 67 638
rect 64 633 67 634
rect 69 638 72 639
rect 84 638 87 639
rect 69 634 70 638
rect 86 634 87 638
rect 69 633 72 634
rect 84 633 87 634
rect 89 638 92 639
rect 89 634 90 638
rect 184 651 187 652
rect 186 647 187 651
rect 184 646 187 647
rect 189 651 192 652
rect 204 651 207 652
rect 189 647 190 651
rect 206 647 207 651
rect 189 646 192 647
rect 204 646 207 647
rect 209 651 212 652
rect 209 647 210 651
rect 209 646 212 647
rect 89 633 92 634
rect 13 624 14 626
rect 18 624 19 626
rect 13 623 19 624
rect 13 620 19 621
rect 13 618 14 620
rect 18 618 19 620
rect 13 604 14 606
rect 18 604 19 606
rect 13 603 19 604
rect 244 638 247 639
rect 246 634 247 638
rect 244 633 247 634
rect 249 638 252 639
rect 264 638 267 639
rect 249 634 250 638
rect 266 634 267 638
rect 249 633 252 634
rect 264 633 267 634
rect 269 638 272 639
rect 269 634 270 638
rect 364 651 367 652
rect 366 647 367 651
rect 364 646 367 647
rect 369 651 372 652
rect 384 651 387 652
rect 369 647 370 651
rect 386 647 387 651
rect 369 646 372 647
rect 384 646 387 647
rect 389 651 392 652
rect 389 647 390 651
rect 389 646 392 647
rect 269 633 272 634
rect 126 612 129 613
rect 128 608 129 612
rect 126 607 129 608
rect 131 612 134 613
rect 146 612 149 613
rect 131 608 132 612
rect 148 608 149 612
rect 131 607 134 608
rect 146 607 149 608
rect 151 612 154 613
rect 597 640 600 641
rect 599 636 600 640
rect 597 635 600 636
rect 602 640 605 641
rect 617 640 620 641
rect 602 636 603 640
rect 619 636 620 640
rect 602 635 605 636
rect 617 635 620 636
rect 622 640 625 641
rect 622 636 623 640
rect 717 653 720 654
rect 719 649 720 653
rect 717 648 720 649
rect 722 653 725 654
rect 737 653 740 654
rect 722 649 723 653
rect 739 649 740 653
rect 722 648 725 649
rect 737 648 740 649
rect 742 653 745 654
rect 742 649 743 653
rect 742 648 745 649
rect 622 635 625 636
rect 151 608 152 612
rect 306 612 309 613
rect 151 607 154 608
rect 308 608 309 612
rect 306 607 309 608
rect 311 612 314 613
rect 326 612 329 613
rect 311 608 312 612
rect 328 608 329 612
rect 311 607 314 608
rect 326 607 329 608
rect 331 612 334 613
rect 777 640 780 641
rect 779 636 780 640
rect 777 635 780 636
rect 782 640 785 641
rect 797 640 800 641
rect 782 636 783 640
rect 799 636 800 640
rect 782 635 785 636
rect 797 635 800 636
rect 802 640 805 641
rect 802 636 803 640
rect 897 653 900 654
rect 899 649 900 653
rect 897 648 900 649
rect 902 653 905 654
rect 917 653 920 654
rect 902 649 903 653
rect 919 649 920 653
rect 902 648 905 649
rect 917 648 920 649
rect 922 653 925 654
rect 922 649 923 653
rect 922 648 925 649
rect 802 635 805 636
rect 407 614 410 615
rect 331 608 332 612
rect 409 610 410 614
rect 407 609 410 610
rect 412 609 426 615
rect 428 614 432 615
rect 441 614 446 615
rect 428 610 429 614
rect 444 610 446 614
rect 428 609 432 610
rect 441 609 446 610
rect 448 614 453 615
rect 448 610 450 614
rect 659 614 662 615
rect 661 610 662 614
rect 448 609 453 610
rect 659 609 662 610
rect 664 614 667 615
rect 679 614 682 615
rect 664 610 665 614
rect 681 610 682 614
rect 664 609 667 610
rect 679 609 682 610
rect 684 614 687 615
rect 684 610 685 614
rect 839 614 842 615
rect 684 609 687 610
rect 841 610 842 614
rect 839 609 842 610
rect 844 614 847 615
rect 859 614 862 615
rect 844 610 845 614
rect 861 610 862 614
rect 844 609 847 610
rect 859 609 862 610
rect 864 614 867 615
rect 939 616 942 617
rect 864 610 865 614
rect 941 612 942 616
rect 939 611 942 612
rect 944 611 958 617
rect 960 616 964 617
rect 973 616 978 617
rect 960 612 961 616
rect 976 612 978 616
rect 960 611 964 612
rect 973 611 978 612
rect 980 616 985 617
rect 980 612 982 616
rect 980 611 985 612
rect 864 609 867 610
rect 331 607 334 608
rect 13 600 19 601
rect 13 598 14 600
rect 18 598 19 600
rect 197 606 200 607
rect 199 602 200 606
rect 197 601 200 602
rect 202 606 206 607
rect 202 602 203 606
rect 202 601 206 602
rect 377 606 380 607
rect 379 602 380 606
rect 377 601 380 602
rect 382 606 386 607
rect 382 602 383 606
rect 382 601 386 602
rect 730 608 733 609
rect 732 604 733 608
rect 730 603 733 604
rect 735 608 739 609
rect 735 604 736 608
rect 735 603 739 604
rect 910 608 913 609
rect 912 604 913 608
rect 910 603 913 604
rect 915 608 919 609
rect 915 604 916 608
rect 915 603 919 604
rect 13 554 14 556
rect 18 554 19 556
rect 13 552 19 554
rect 13 549 19 550
rect 13 546 14 549
rect 18 546 19 549
rect 13 537 14 539
rect 18 537 19 539
rect 13 536 19 537
rect 13 533 19 534
rect 13 531 14 533
rect 18 531 19 533
rect 13 517 14 519
rect 18 517 19 519
rect 13 516 19 517
rect 13 513 19 514
rect 13 511 14 513
rect 18 511 19 513
rect 317 506 320 507
rect 319 502 320 506
rect 317 501 320 502
rect 322 506 325 507
rect 337 506 340 507
rect 322 502 323 506
rect 339 502 340 506
rect 322 501 325 502
rect 337 501 340 502
rect 342 506 345 507
rect 497 506 500 507
rect 342 502 343 506
rect 499 502 500 506
rect 342 501 345 502
rect 497 501 500 502
rect 502 506 505 507
rect 517 506 520 507
rect 502 502 503 506
rect 519 502 520 506
rect 502 501 505 502
rect 517 501 520 502
rect 522 506 525 507
rect 522 502 523 506
rect 522 501 525 502
rect 255 483 258 484
rect 257 479 258 483
rect 255 478 258 479
rect 260 483 263 484
rect 275 483 278 484
rect 260 479 261 483
rect 277 479 278 483
rect 260 478 263 479
rect 275 478 278 479
rect 280 483 283 484
rect 280 479 281 483
rect 375 496 378 497
rect 377 492 378 496
rect 375 491 378 492
rect 380 496 383 497
rect 395 496 398 497
rect 380 492 381 496
rect 397 492 398 496
rect 380 491 383 492
rect 395 491 398 492
rect 400 496 403 497
rect 400 492 401 496
rect 400 491 403 492
rect 280 478 283 479
rect 14 466 15 468
rect 19 466 20 468
rect 14 464 20 466
rect 14 461 20 462
rect 14 458 15 461
rect 19 458 20 461
rect 435 483 438 484
rect 437 479 438 483
rect 435 478 438 479
rect 440 483 443 484
rect 455 483 458 484
rect 440 479 441 483
rect 457 479 458 483
rect 440 478 443 479
rect 455 478 458 479
rect 460 483 463 484
rect 460 479 461 483
rect 555 496 558 497
rect 557 492 558 496
rect 555 491 558 492
rect 560 496 563 497
rect 575 496 578 497
rect 560 492 561 496
rect 577 492 578 496
rect 560 491 563 492
rect 575 491 578 492
rect 580 496 583 497
rect 580 492 581 496
rect 580 491 583 492
rect 460 478 463 479
rect 317 457 320 458
rect 319 453 320 457
rect 14 449 15 451
rect 19 449 20 451
rect 317 452 320 453
rect 322 457 325 458
rect 337 457 340 458
rect 322 453 323 457
rect 339 453 340 457
rect 322 452 325 453
rect 337 452 340 453
rect 342 457 345 458
rect 342 453 343 457
rect 497 457 500 458
rect 342 452 345 453
rect 499 453 500 457
rect 497 452 500 453
rect 502 457 505 458
rect 517 457 520 458
rect 502 453 503 457
rect 519 453 520 457
rect 502 452 505 453
rect 517 452 520 453
rect 522 457 525 458
rect 597 459 600 460
rect 522 453 523 457
rect 599 455 600 459
rect 597 454 600 455
rect 602 454 616 460
rect 618 459 622 460
rect 631 459 636 460
rect 618 455 619 459
rect 634 455 636 459
rect 618 454 622 455
rect 631 454 636 455
rect 638 459 643 460
rect 638 455 640 459
rect 638 454 643 455
rect 522 452 525 453
rect 14 448 20 449
rect 14 445 20 446
rect 14 443 15 445
rect 19 443 20 445
rect 14 429 15 431
rect 19 429 20 431
rect 14 428 20 429
rect 388 451 391 452
rect 390 447 391 451
rect 388 446 391 447
rect 393 451 397 452
rect 393 447 394 451
rect 393 446 397 447
rect 568 451 571 452
rect 570 447 571 451
rect 568 446 571 447
rect 573 451 577 452
rect 573 447 574 451
rect 573 446 577 447
rect 14 425 20 426
rect 14 423 15 425
rect 19 423 20 425
rect 147 405 150 406
rect 149 401 150 405
rect 147 400 150 401
rect 152 405 155 406
rect 167 405 170 406
rect 152 401 153 405
rect 169 401 170 405
rect 152 400 155 401
rect 167 400 170 401
rect 172 405 175 406
rect 172 401 173 405
rect 172 400 175 401
rect 15 385 16 387
rect 20 385 21 387
rect 15 383 21 385
rect 15 380 21 381
rect 15 377 16 380
rect 20 377 21 380
rect 85 382 88 383
rect 87 378 88 382
rect 85 377 88 378
rect 90 382 93 383
rect 105 382 108 383
rect 90 378 91 382
rect 107 378 108 382
rect 90 377 93 378
rect 105 377 108 378
rect 110 382 113 383
rect 110 378 111 382
rect 205 395 208 396
rect 207 391 208 395
rect 205 390 208 391
rect 210 395 213 396
rect 225 395 228 396
rect 210 391 211 395
rect 227 391 228 395
rect 210 390 213 391
rect 225 390 228 391
rect 230 395 233 396
rect 230 391 231 395
rect 230 390 233 391
rect 110 377 113 378
rect 15 368 16 370
rect 20 368 21 370
rect 15 367 21 368
rect 15 364 21 365
rect 15 362 16 364
rect 20 362 21 364
rect 15 348 16 350
rect 20 348 21 350
rect 15 347 21 348
rect 564 371 567 372
rect 566 367 567 371
rect 564 366 567 367
rect 569 371 572 372
rect 584 371 587 372
rect 569 367 570 371
rect 586 367 587 371
rect 569 366 572 367
rect 584 366 587 367
rect 589 371 592 372
rect 744 371 747 372
rect 589 367 590 371
rect 746 367 747 371
rect 589 366 592 367
rect 744 366 747 367
rect 749 371 752 372
rect 764 371 767 372
rect 749 367 750 371
rect 766 367 767 371
rect 749 366 752 367
rect 764 366 767 367
rect 769 371 772 372
rect 769 367 770 371
rect 769 366 772 367
rect 147 356 150 357
rect 149 352 150 356
rect 147 351 150 352
rect 152 356 155 357
rect 167 356 170 357
rect 152 352 153 356
rect 169 352 170 356
rect 152 351 155 352
rect 167 351 170 352
rect 172 356 175 357
rect 172 352 173 356
rect 172 351 175 352
rect 15 344 21 345
rect 15 342 16 344
rect 20 342 21 344
rect 218 350 221 351
rect 220 346 221 350
rect 218 345 221 346
rect 223 350 227 351
rect 223 346 224 350
rect 502 348 505 349
rect 223 345 227 346
rect 504 344 505 348
rect 502 343 505 344
rect 507 348 510 349
rect 522 348 525 349
rect 507 344 508 348
rect 524 344 525 348
rect 507 343 510 344
rect 522 343 525 344
rect 527 348 530 349
rect 527 344 528 348
rect 622 361 625 362
rect 624 357 625 361
rect 622 356 625 357
rect 627 361 630 362
rect 642 361 645 362
rect 627 357 628 361
rect 644 357 645 361
rect 627 356 630 357
rect 642 356 645 357
rect 647 361 650 362
rect 647 357 648 361
rect 647 356 650 357
rect 527 343 530 344
rect 682 348 685 349
rect 684 344 685 348
rect 682 343 685 344
rect 687 348 690 349
rect 702 348 705 349
rect 687 344 688 348
rect 704 344 705 348
rect 687 343 690 344
rect 702 343 705 344
rect 707 348 710 349
rect 707 344 708 348
rect 802 361 805 362
rect 804 357 805 361
rect 802 356 805 357
rect 807 361 810 362
rect 822 361 825 362
rect 807 357 808 361
rect 824 357 825 361
rect 807 356 810 357
rect 822 356 825 357
rect 827 361 830 362
rect 827 357 828 361
rect 827 356 830 357
rect 707 343 710 344
rect 564 322 567 323
rect 566 318 567 322
rect 564 317 567 318
rect 569 322 572 323
rect 584 322 587 323
rect 569 318 570 322
rect 586 318 587 322
rect 569 317 572 318
rect 584 317 587 318
rect 589 322 592 323
rect 589 318 590 322
rect 744 322 747 323
rect 589 317 592 318
rect 746 318 747 322
rect 744 317 747 318
rect 749 322 752 323
rect 764 322 767 323
rect 749 318 750 322
rect 766 318 767 322
rect 749 317 752 318
rect 764 317 767 318
rect 769 322 772 323
rect 844 324 847 325
rect 769 318 770 322
rect 846 320 847 324
rect 844 319 847 320
rect 849 319 863 325
rect 865 324 869 325
rect 878 324 883 325
rect 865 320 866 324
rect 881 320 883 324
rect 865 319 869 320
rect 878 319 883 320
rect 885 324 890 325
rect 885 320 887 324
rect 885 319 890 320
rect 769 317 772 318
rect 15 301 16 303
rect 20 301 21 303
rect 15 299 21 301
rect 15 296 21 297
rect 15 293 16 296
rect 20 293 21 296
rect 635 316 638 317
rect 637 312 638 316
rect 635 311 638 312
rect 640 316 644 317
rect 640 312 641 316
rect 640 311 644 312
rect 815 316 818 317
rect 817 312 818 316
rect 815 311 818 312
rect 820 316 824 317
rect 820 312 821 316
rect 820 311 824 312
rect 15 284 16 286
rect 20 284 21 286
rect 15 283 21 284
rect 15 280 21 281
rect 15 278 16 280
rect 20 278 21 280
rect 15 264 16 266
rect 20 264 21 266
rect 15 263 21 264
rect 15 260 21 261
rect 15 258 16 260
rect 20 258 21 260
rect 164 219 167 220
rect 15 214 16 216
rect 20 214 21 216
rect 15 212 21 214
rect 166 215 167 219
rect 164 214 167 215
rect 169 219 172 220
rect 184 219 187 220
rect 169 215 170 219
rect 186 215 187 219
rect 169 214 172 215
rect 184 214 187 215
rect 189 219 192 220
rect 344 219 347 220
rect 189 215 190 219
rect 346 215 347 219
rect 189 214 192 215
rect 344 214 347 215
rect 349 219 352 220
rect 364 219 367 220
rect 349 215 350 219
rect 366 215 367 219
rect 349 214 352 215
rect 364 214 367 215
rect 369 219 372 220
rect 369 215 370 219
rect 369 214 372 215
rect 15 209 21 210
rect 15 206 16 209
rect 20 206 21 209
rect 15 197 16 199
rect 20 197 21 199
rect 15 196 21 197
rect 102 196 105 197
rect 15 193 21 194
rect 15 191 16 193
rect 20 191 21 193
rect 15 177 16 179
rect 20 177 21 179
rect 15 176 21 177
rect 104 192 105 196
rect 102 191 105 192
rect 107 196 110 197
rect 122 196 125 197
rect 107 192 108 196
rect 124 192 125 196
rect 107 191 110 192
rect 122 191 125 192
rect 127 196 130 197
rect 127 192 128 196
rect 222 209 225 210
rect 224 205 225 209
rect 222 204 225 205
rect 227 209 230 210
rect 242 209 245 210
rect 227 205 228 209
rect 244 205 245 209
rect 227 204 230 205
rect 242 204 245 205
rect 247 209 250 210
rect 247 205 248 209
rect 247 204 250 205
rect 127 191 130 192
rect 15 173 21 174
rect 15 171 16 173
rect 20 171 21 173
rect 282 196 285 197
rect 284 192 285 196
rect 282 191 285 192
rect 287 196 290 197
rect 302 196 305 197
rect 287 192 288 196
rect 304 192 305 196
rect 287 191 290 192
rect 302 191 305 192
rect 307 196 310 197
rect 307 192 308 196
rect 402 209 405 210
rect 404 205 405 209
rect 402 204 405 205
rect 407 209 410 210
rect 422 209 425 210
rect 407 205 408 209
rect 424 205 425 209
rect 407 204 410 205
rect 422 204 425 205
rect 427 209 430 210
rect 427 205 428 209
rect 427 204 430 205
rect 307 191 310 192
rect 164 170 167 171
rect 166 166 167 170
rect 164 165 167 166
rect 169 170 172 171
rect 184 170 187 171
rect 169 166 170 170
rect 186 166 187 170
rect 169 165 172 166
rect 184 165 187 166
rect 189 170 192 171
rect 189 166 190 170
rect 344 170 347 171
rect 189 165 192 166
rect 346 166 347 170
rect 344 165 347 166
rect 349 170 352 171
rect 364 170 367 171
rect 349 166 350 170
rect 366 166 367 170
rect 349 165 352 166
rect 364 165 367 166
rect 369 170 372 171
rect 444 172 447 173
rect 369 166 370 170
rect 446 168 447 172
rect 444 167 447 168
rect 449 167 463 173
rect 465 172 469 173
rect 478 172 483 173
rect 465 168 466 172
rect 481 168 483 172
rect 465 167 469 168
rect 478 167 483 168
rect 485 172 490 173
rect 587 172 590 173
rect 485 168 487 172
rect 589 168 590 172
rect 485 167 490 168
rect 587 167 590 168
rect 592 172 595 173
rect 607 172 610 173
rect 592 168 593 172
rect 609 168 610 172
rect 592 167 595 168
rect 607 167 610 168
rect 612 172 615 173
rect 767 172 770 173
rect 612 168 613 172
rect 769 168 770 172
rect 612 167 615 168
rect 767 167 770 168
rect 772 172 775 173
rect 787 172 790 173
rect 772 168 773 172
rect 789 168 790 172
rect 772 167 775 168
rect 787 167 790 168
rect 792 172 795 173
rect 792 168 793 172
rect 792 167 795 168
rect 369 165 372 166
rect 235 164 238 165
rect 237 160 238 164
rect 235 159 238 160
rect 240 164 244 165
rect 240 160 241 164
rect 240 159 244 160
rect 415 164 418 165
rect 417 160 418 164
rect 415 159 418 160
rect 420 164 424 165
rect 420 160 421 164
rect 420 159 424 160
rect 525 149 528 150
rect 527 145 528 149
rect 525 144 528 145
rect 530 149 533 150
rect 545 149 548 150
rect 530 145 531 149
rect 547 145 548 149
rect 530 144 533 145
rect 545 144 548 145
rect 550 149 553 150
rect 550 145 551 149
rect 645 162 648 163
rect 647 158 648 162
rect 645 157 648 158
rect 650 162 653 163
rect 665 162 668 163
rect 650 158 651 162
rect 667 158 668 162
rect 650 157 653 158
rect 665 157 668 158
rect 670 162 673 163
rect 670 158 671 162
rect 670 157 673 158
rect 550 144 553 145
rect 16 126 17 128
rect 21 126 22 128
rect 16 124 22 126
rect 705 149 708 150
rect 707 145 708 149
rect 705 144 708 145
rect 710 149 713 150
rect 725 149 728 150
rect 710 145 711 149
rect 727 145 728 149
rect 710 144 713 145
rect 725 144 728 145
rect 730 149 733 150
rect 730 145 731 149
rect 825 162 828 163
rect 827 158 828 162
rect 825 157 828 158
rect 830 162 833 163
rect 845 162 848 163
rect 830 158 831 162
rect 847 158 848 162
rect 830 157 833 158
rect 845 157 848 158
rect 850 162 853 163
rect 850 158 851 162
rect 850 157 853 158
rect 730 144 733 145
rect 16 121 22 122
rect 16 118 17 121
rect 21 118 22 121
rect 587 123 590 124
rect 589 119 590 123
rect 587 118 590 119
rect 592 123 595 124
rect 607 123 610 124
rect 592 119 593 123
rect 609 119 610 123
rect 592 118 595 119
rect 607 118 610 119
rect 612 123 615 124
rect 612 119 613 123
rect 767 123 770 124
rect 612 118 615 119
rect 769 119 770 123
rect 767 118 770 119
rect 772 123 775 124
rect 787 123 790 124
rect 772 119 773 123
rect 789 119 790 123
rect 772 118 775 119
rect 787 118 790 119
rect 792 123 795 124
rect 867 125 870 126
rect 792 119 793 123
rect 869 121 870 125
rect 867 120 870 121
rect 872 120 886 126
rect 888 125 892 126
rect 901 125 906 126
rect 888 121 889 125
rect 904 121 906 125
rect 888 120 892 121
rect 901 120 906 121
rect 908 125 913 126
rect 908 121 910 125
rect 908 120 913 121
rect 792 118 795 119
rect 16 109 17 111
rect 21 109 22 111
rect 16 108 22 109
rect 16 105 22 106
rect 16 103 17 105
rect 21 103 22 105
rect 16 89 17 91
rect 21 89 22 91
rect 16 88 22 89
rect 658 117 661 118
rect 660 113 661 117
rect 658 112 661 113
rect 663 117 667 118
rect 663 113 664 117
rect 663 112 667 113
rect 838 117 841 118
rect 840 113 841 117
rect 838 112 841 113
rect 843 117 847 118
rect 843 113 844 117
rect 843 112 847 113
rect 16 85 22 86
rect 16 83 17 85
rect 21 83 22 85
rect 17 45 18 47
rect 22 45 23 47
rect 17 43 23 45
rect 17 40 23 41
rect 17 37 18 40
rect 22 37 23 40
rect 17 28 18 30
rect 22 28 23 30
rect 17 27 23 28
rect 17 24 23 25
rect 17 22 18 24
rect 22 22 23 24
rect 17 8 18 10
rect 22 8 23 10
rect 17 7 23 8
rect 17 4 23 5
rect 17 2 18 4
rect 22 2 23 4
<< metal1 >>
rect 14 1321 31 1324
rect 4 1312 10 1315
rect 1 1300 4 1312
rect 17 1308 20 1314
rect 35 1312 39 1315
rect 14 1305 31 1308
rect 4 1296 10 1299
rect 1 1280 4 1296
rect 17 1288 20 1305
rect 14 1285 20 1288
rect 4 1277 10 1280
rect 40 1280 43 1311
rect 35 1276 39 1279
rect 0 1263 3 1276
rect 0 1229 3 1259
rect 26 1237 29 1242
rect 14 1234 31 1237
rect 4 1225 10 1228
rect 1 1213 4 1225
rect 17 1221 20 1227
rect 40 1228 43 1276
rect 91 1259 131 1262
rect 135 1259 139 1262
rect 143 1259 159 1262
rect 163 1259 197 1262
rect 201 1260 315 1262
rect 319 1260 359 1263
rect 363 1260 367 1263
rect 371 1260 387 1263
rect 391 1260 425 1263
rect 429 1260 464 1263
rect 201 1259 319 1260
rect 140 1253 143 1259
rect 159 1253 162 1259
rect 198 1253 201 1259
rect 201 1249 217 1252
rect 148 1246 151 1249
rect 168 1246 171 1249
rect 60 1243 141 1246
rect 35 1225 39 1228
rect 14 1218 31 1221
rect 4 1209 10 1212
rect 1 1193 4 1209
rect 17 1201 20 1218
rect 14 1198 20 1201
rect 4 1190 10 1193
rect 40 1193 43 1224
rect 71 1223 74 1243
rect 148 1243 171 1246
rect 198 1243 201 1249
rect 217 1243 220 1249
rect 81 1236 87 1239
rect 91 1236 97 1239
rect 78 1230 81 1236
rect 97 1230 100 1236
rect 115 1235 161 1238
rect 168 1236 171 1243
rect 206 1236 209 1239
rect 226 1236 229 1239
rect 86 1223 89 1226
rect 106 1223 109 1226
rect 115 1223 118 1235
rect 168 1233 199 1236
rect 168 1232 171 1233
rect 206 1233 229 1236
rect 139 1224 142 1228
rect 174 1225 219 1228
rect 71 1220 79 1223
rect 86 1220 118 1223
rect 128 1220 139 1223
rect 35 1189 39 1192
rect 1 1141 4 1189
rect 40 1176 43 1189
rect 71 1213 99 1216
rect 71 1190 74 1213
rect 106 1209 109 1220
rect 77 1197 80 1205
rect 115 1198 118 1220
rect 135 1210 139 1213
rect 143 1210 159 1213
rect 140 1204 143 1210
rect 159 1204 162 1210
rect 148 1197 151 1200
rect 168 1197 171 1200
rect 174 1197 177 1225
rect 226 1222 229 1233
rect 119 1194 141 1197
rect 148 1194 177 1197
rect 71 1187 161 1190
rect 27 1149 30 1154
rect 15 1146 32 1149
rect 5 1137 11 1140
rect 2 1125 5 1137
rect 18 1133 21 1139
rect 40 1140 43 1172
rect 71 1160 74 1187
rect 168 1183 171 1194
rect 139 1175 142 1179
rect 197 1175 200 1218
rect 210 1204 221 1205
rect 233 1207 236 1259
rect 368 1254 371 1260
rect 387 1254 390 1260
rect 426 1254 429 1260
rect 429 1250 445 1253
rect 376 1247 379 1250
rect 396 1247 399 1250
rect 225 1204 236 1207
rect 258 1244 369 1247
rect 210 1202 224 1204
rect 210 1198 213 1202
rect 222 1194 224 1198
rect 221 1192 224 1194
rect 258 1192 261 1244
rect 299 1224 302 1244
rect 376 1244 399 1247
rect 426 1244 429 1250
rect 445 1244 448 1250
rect 309 1237 315 1240
rect 319 1237 325 1240
rect 306 1231 309 1237
rect 325 1231 328 1237
rect 343 1236 389 1239
rect 396 1237 399 1244
rect 434 1237 437 1240
rect 454 1237 457 1240
rect 314 1224 317 1227
rect 334 1224 337 1227
rect 343 1224 346 1236
rect 396 1234 427 1237
rect 396 1233 399 1234
rect 434 1234 457 1237
rect 367 1225 370 1229
rect 402 1226 447 1229
rect 299 1221 307 1224
rect 314 1221 346 1224
rect 356 1221 367 1224
rect 299 1214 327 1217
rect 299 1192 302 1214
rect 334 1210 337 1221
rect 305 1198 308 1206
rect 343 1199 346 1221
rect 363 1211 367 1214
rect 371 1211 387 1214
rect 368 1205 371 1211
rect 387 1205 390 1211
rect 376 1198 379 1201
rect 396 1198 399 1201
rect 402 1198 405 1226
rect 454 1223 457 1234
rect 347 1195 369 1198
rect 376 1195 405 1198
rect 207 1186 213 1189
rect 221 1189 261 1192
rect 221 1182 224 1189
rect 301 1191 302 1192
rect 301 1188 389 1191
rect 396 1184 399 1195
rect 223 1178 224 1182
rect 209 1175 212 1178
rect 367 1176 370 1180
rect 425 1176 428 1219
rect 438 1205 449 1206
rect 461 1208 464 1260
rect 453 1205 464 1208
rect 438 1203 452 1205
rect 438 1199 441 1203
rect 450 1195 452 1199
rect 435 1187 441 1190
rect 449 1190 452 1195
rect 449 1185 451 1190
rect 449 1183 452 1185
rect 451 1179 452 1183
rect 437 1176 440 1179
rect 81 1172 99 1175
rect 103 1172 125 1175
rect 129 1172 139 1175
rect 143 1172 167 1175
rect 171 1172 196 1175
rect 200 1174 305 1175
rect 200 1172 219 1174
rect 223 1172 305 1174
rect 309 1173 327 1176
rect 331 1173 353 1176
rect 357 1173 367 1176
rect 371 1173 395 1176
rect 399 1173 424 1176
rect 428 1175 450 1176
rect 428 1173 447 1175
rect 36 1137 40 1140
rect 15 1130 32 1133
rect 5 1121 11 1124
rect 2 1105 5 1121
rect 18 1113 21 1130
rect 15 1110 21 1113
rect 5 1102 11 1105
rect 41 1105 44 1136
rect 36 1101 40 1104
rect 2 1060 5 1101
rect 28 1068 31 1073
rect 16 1065 33 1068
rect 6 1056 12 1059
rect 3 1044 6 1056
rect 19 1052 22 1058
rect 41 1059 44 1101
rect 37 1056 41 1059
rect 16 1049 33 1052
rect 6 1040 12 1043
rect 3 1024 6 1040
rect 19 1032 22 1049
rect 16 1029 22 1032
rect 6 1021 12 1024
rect 42 1024 45 1055
rect 37 1020 41 1023
rect 3 1009 6 1020
rect 3 976 6 1005
rect 28 984 31 989
rect 16 981 33 984
rect 6 972 12 975
rect 3 960 6 972
rect 19 968 22 974
rect 42 975 45 1020
rect 78 1005 118 1008
rect 122 1005 126 1008
rect 130 1005 146 1008
rect 150 1005 184 1008
rect 188 1005 254 1008
rect 258 1005 298 1008
rect 302 1005 306 1008
rect 310 1005 326 1008
rect 330 1005 364 1008
rect 368 1005 404 1008
rect 127 999 130 1005
rect 146 999 149 1005
rect 185 999 188 1005
rect 188 995 204 998
rect 37 972 41 975
rect 16 965 33 968
rect 6 956 12 959
rect 3 940 6 956
rect 19 948 22 965
rect 16 945 22 948
rect 6 937 12 940
rect 42 940 45 971
rect 135 992 138 995
rect 155 992 158 995
rect 62 989 128 992
rect 58 969 61 989
rect 135 989 158 992
rect 185 989 188 995
rect 204 989 207 995
rect 68 982 74 985
rect 78 982 84 985
rect 65 976 68 982
rect 84 976 87 982
rect 102 981 148 984
rect 155 982 158 989
rect 193 982 196 985
rect 213 982 216 985
rect 73 969 76 972
rect 93 969 96 972
rect 102 969 105 981
rect 155 979 186 982
rect 155 978 158 979
rect 193 979 216 982
rect 213 978 216 979
rect 126 970 129 974
rect 161 971 206 974
rect 213 974 214 978
rect 58 966 66 969
rect 73 966 105 969
rect 115 966 126 969
rect 37 936 41 939
rect 58 959 86 962
rect 58 937 61 959
rect 93 955 96 966
rect 64 943 67 951
rect 102 944 105 966
rect 122 956 126 959
rect 130 956 146 959
rect 127 950 130 956
rect 146 950 149 956
rect 135 943 138 946
rect 155 943 158 946
rect 161 943 164 971
rect 213 968 216 974
rect 106 940 128 943
rect 135 940 164 943
rect 3 889 6 936
rect 41 921 44 936
rect 60 936 61 937
rect 60 933 148 936
rect 155 929 158 940
rect 126 921 129 925
rect 184 921 187 964
rect 197 950 208 951
rect 222 953 225 1005
rect 307 999 310 1005
rect 326 999 329 1005
rect 365 999 368 1005
rect 368 995 384 998
rect 315 992 318 995
rect 335 992 338 995
rect 242 989 308 992
rect 238 969 241 989
rect 315 989 338 992
rect 365 989 368 995
rect 384 989 387 995
rect 248 982 254 985
rect 258 982 264 985
rect 245 976 248 982
rect 264 976 267 982
rect 282 981 328 984
rect 335 982 338 989
rect 373 982 376 985
rect 393 982 396 985
rect 253 969 256 972
rect 273 969 276 972
rect 282 969 285 981
rect 335 979 366 982
rect 335 978 338 979
rect 373 980 396 982
rect 373 979 394 980
rect 393 976 394 979
rect 306 970 309 974
rect 341 971 386 974
rect 238 966 246 969
rect 253 966 285 969
rect 295 966 306 969
rect 212 950 225 953
rect 238 959 266 962
rect 238 951 241 959
rect 273 955 276 966
rect 197 948 211 950
rect 197 944 200 948
rect 240 946 241 951
rect 209 940 211 944
rect 194 932 200 935
rect 208 935 211 940
rect 238 936 241 946
rect 244 943 247 951
rect 282 944 285 966
rect 302 956 306 959
rect 310 956 326 959
rect 307 950 310 956
rect 326 950 329 956
rect 315 943 318 946
rect 335 943 338 946
rect 341 943 344 971
rect 393 968 396 976
rect 286 940 308 943
rect 315 940 344 943
rect 208 931 209 935
rect 238 933 328 936
rect 208 928 211 931
rect 335 929 338 940
rect 210 924 211 928
rect 196 921 199 924
rect 306 921 309 925
rect 364 921 367 964
rect 401 961 404 1005
rect 436 1002 569 1005
rect 573 1002 613 1005
rect 617 1002 621 1005
rect 625 1002 641 1005
rect 645 1002 679 1005
rect 683 1002 718 1005
rect 436 961 439 1002
rect 622 996 625 1002
rect 641 996 644 1002
rect 680 996 683 1002
rect 683 992 699 995
rect 553 986 560 989
rect 630 989 633 992
rect 650 989 653 992
rect 565 986 623 989
rect 553 966 556 986
rect 630 986 653 989
rect 680 986 683 992
rect 699 986 702 992
rect 563 979 569 982
rect 573 979 579 982
rect 560 973 563 979
rect 579 973 582 979
rect 597 978 643 981
rect 650 979 653 986
rect 688 979 691 982
rect 708 979 711 982
rect 568 966 571 969
rect 588 966 591 969
rect 597 966 600 978
rect 650 976 681 979
rect 650 975 653 976
rect 688 976 711 979
rect 621 967 624 971
rect 656 968 701 971
rect 553 963 561 966
rect 568 963 600 966
rect 610 963 621 966
rect 401 958 407 961
rect 377 950 388 951
rect 401 953 404 958
rect 392 950 404 953
rect 411 958 442 961
rect 407 952 410 957
rect 442 952 445 957
rect 552 956 581 959
rect 377 948 391 950
rect 377 944 380 948
rect 389 943 391 944
rect 389 940 425 943
rect 374 932 380 935
rect 388 928 391 940
rect 401 931 409 934
rect 432 934 435 948
rect 453 937 456 948
rect 416 931 446 934
rect 453 933 474 937
rect 552 934 555 956
rect 588 952 591 963
rect 559 940 562 948
rect 597 941 600 963
rect 617 953 621 956
rect 625 953 641 956
rect 622 947 625 953
rect 641 947 644 953
rect 630 940 633 943
rect 650 940 653 943
rect 656 940 659 968
rect 708 965 711 976
rect 601 937 623 940
rect 630 937 659 940
rect 416 928 419 931
rect 432 928 435 931
rect 453 928 456 933
rect 390 924 391 928
rect 376 921 379 924
rect 407 921 410 924
rect 423 921 426 924
rect 443 921 446 924
rect 41 918 64 921
rect 29 897 32 902
rect 16 894 33 897
rect 6 885 12 888
rect 3 873 6 885
rect 19 881 22 887
rect 41 888 44 918
rect 68 918 86 921
rect 90 918 112 921
rect 116 918 126 921
rect 130 918 154 921
rect 158 918 183 921
rect 187 920 244 921
rect 187 918 206 920
rect 210 918 244 920
rect 248 918 266 921
rect 270 918 292 921
rect 296 918 306 921
rect 310 918 334 921
rect 338 918 363 921
rect 367 920 446 921
rect 367 918 386 920
rect 390 918 419 920
rect 423 918 446 920
rect 224 906 397 909
rect 430 895 433 918
rect 471 906 474 933
rect 555 930 643 933
rect 650 926 653 937
rect 621 918 624 922
rect 679 918 682 961
rect 692 947 703 948
rect 715 950 718 1002
rect 707 947 718 950
rect 692 945 706 947
rect 692 941 695 945
rect 704 937 706 941
rect 689 929 695 932
rect 703 929 706 937
rect 703 926 820 929
rect 703 925 706 926
rect 705 921 706 925
rect 691 918 694 921
rect 543 915 559 918
rect 543 895 546 915
rect 563 915 581 918
rect 585 915 607 918
rect 611 915 621 918
rect 625 915 649 918
rect 653 915 678 918
rect 682 917 704 918
rect 682 915 701 917
rect 430 892 546 895
rect 37 885 41 888
rect 16 878 33 881
rect 6 869 12 872
rect 3 853 6 869
rect 19 861 22 878
rect 16 858 22 861
rect 6 850 12 853
rect 42 853 45 884
rect 37 849 41 852
rect 3 838 6 849
rect 3 801 6 833
rect 29 809 32 814
rect 17 806 34 809
rect 7 797 13 800
rect 4 785 7 797
rect 20 793 23 799
rect 42 800 45 849
rect 281 834 321 837
rect 325 834 329 837
rect 333 834 349 837
rect 353 834 387 837
rect 391 834 457 837
rect 461 834 501 837
rect 505 834 509 837
rect 513 834 529 837
rect 533 834 567 837
rect 571 834 606 837
rect 330 828 333 834
rect 349 828 352 834
rect 388 828 391 834
rect 391 824 407 827
rect 338 821 341 824
rect 358 821 361 824
rect 261 818 331 821
rect 38 797 42 800
rect 17 790 34 793
rect 7 781 13 784
rect 4 765 7 781
rect 20 773 23 790
rect 17 770 23 773
rect 7 762 13 765
rect 43 765 46 796
rect 261 798 264 818
rect 338 818 361 821
rect 388 818 391 824
rect 407 818 410 824
rect 271 811 277 814
rect 281 811 287 814
rect 268 805 271 811
rect 287 805 290 811
rect 305 810 351 813
rect 358 811 361 818
rect 396 811 399 814
rect 416 811 419 814
rect 276 798 279 801
rect 296 798 299 801
rect 305 798 308 810
rect 358 808 389 811
rect 358 807 361 808
rect 396 808 419 811
rect 416 807 419 808
rect 329 799 332 803
rect 364 800 409 803
rect 416 803 417 807
rect 261 795 269 798
rect 276 795 308 798
rect 318 795 329 798
rect 261 788 289 791
rect 261 766 264 788
rect 296 784 299 795
rect 267 772 270 780
rect 305 773 308 795
rect 325 785 329 788
rect 333 785 349 788
rect 330 779 333 785
rect 349 779 352 785
rect 338 772 341 775
rect 358 772 361 775
rect 364 772 367 800
rect 416 797 419 803
rect 309 769 331 772
rect 338 769 367 772
rect 38 761 42 764
rect 263 765 264 766
rect 263 762 351 765
rect 4 720 7 761
rect 43 750 46 761
rect 358 758 361 769
rect 329 750 332 754
rect 387 750 390 793
rect 400 779 411 780
rect 425 782 428 834
rect 510 828 513 834
rect 529 828 532 834
rect 568 828 571 834
rect 571 824 587 827
rect 518 821 521 824
rect 538 821 541 824
rect 445 818 511 821
rect 441 798 444 818
rect 518 818 541 821
rect 568 818 571 824
rect 587 818 590 824
rect 451 811 457 814
rect 461 811 467 814
rect 448 805 451 811
rect 467 805 470 811
rect 485 810 531 813
rect 538 811 541 818
rect 576 811 579 814
rect 596 811 599 814
rect 456 798 459 801
rect 476 798 479 801
rect 485 798 488 810
rect 538 808 569 811
rect 538 807 541 808
rect 576 810 599 811
rect 576 808 596 810
rect 509 799 512 803
rect 544 800 589 803
rect 441 795 449 798
rect 456 795 488 798
rect 498 795 509 798
rect 415 779 428 782
rect 441 788 469 791
rect 441 780 444 788
rect 476 784 479 795
rect 400 777 414 779
rect 400 773 403 777
rect 443 775 444 780
rect 412 769 414 773
rect 397 761 403 764
rect 411 764 414 769
rect 441 765 444 775
rect 447 772 450 780
rect 485 773 488 795
rect 505 785 509 788
rect 513 785 529 788
rect 510 779 513 785
rect 529 779 532 785
rect 518 772 521 775
rect 538 772 541 775
rect 544 772 547 800
rect 596 797 599 806
rect 489 769 511 772
rect 518 769 547 772
rect 411 760 412 764
rect 441 762 531 765
rect 411 757 414 760
rect 538 758 541 769
rect 413 753 414 757
rect 399 750 402 753
rect 509 750 512 754
rect 567 750 570 793
rect 603 790 606 834
rect 603 787 609 790
rect 580 779 591 780
rect 603 782 606 787
rect 595 779 606 782
rect 613 787 644 790
rect 609 781 612 786
rect 644 781 647 786
rect 580 777 594 779
rect 580 773 583 777
rect 592 772 594 773
rect 592 769 627 772
rect 577 761 583 764
rect 591 757 594 769
rect 604 760 611 763
rect 634 763 637 777
rect 618 760 648 763
rect 655 763 658 777
rect 655 760 667 763
rect 618 757 621 760
rect 634 757 637 760
rect 655 757 658 760
rect 593 753 594 757
rect 579 750 582 753
rect 609 750 612 753
rect 625 750 628 753
rect 645 750 648 753
rect 43 747 267 750
rect 31 728 34 734
rect 18 725 35 728
rect 8 716 14 719
rect 5 704 8 716
rect 21 712 24 718
rect 43 719 46 747
rect 271 747 289 750
rect 293 747 315 750
rect 319 747 329 750
rect 333 747 357 750
rect 361 747 386 750
rect 390 749 447 750
rect 390 747 409 749
rect 413 747 447 749
rect 451 747 469 750
rect 473 747 495 750
rect 499 747 509 750
rect 513 747 537 750
rect 541 747 566 750
rect 570 749 648 750
rect 570 747 589 749
rect 593 747 621 749
rect 625 747 648 749
rect 427 735 600 738
rect 664 734 667 760
rect 640 731 667 734
rect 39 716 43 719
rect 18 709 35 712
rect 8 700 14 703
rect 5 684 8 700
rect 21 692 24 709
rect 18 689 24 692
rect 8 681 14 684
rect 44 684 47 715
rect 39 680 43 683
rect 640 688 643 731
rect 817 695 820 926
rect 5 670 8 680
rect 5 636 8 666
rect 31 644 34 650
rect 18 641 35 644
rect 8 632 14 635
rect 5 620 8 632
rect 21 628 24 634
rect 43 635 46 680
rect 76 667 116 670
rect 120 667 124 670
rect 128 667 144 670
rect 148 667 182 670
rect 186 667 252 670
rect 256 667 296 670
rect 300 667 304 670
rect 308 667 324 670
rect 328 667 362 670
rect 366 667 402 670
rect 125 661 128 667
rect 144 661 147 667
rect 183 661 186 667
rect 186 657 202 660
rect 133 654 136 657
rect 153 654 156 657
rect 59 651 126 654
rect 39 632 43 635
rect 18 625 35 628
rect 8 616 14 619
rect 5 600 8 616
rect 21 608 24 625
rect 18 605 24 608
rect 8 597 14 600
rect 44 600 47 631
rect 56 631 59 651
rect 133 651 156 654
rect 183 651 186 657
rect 202 651 205 657
rect 66 644 72 647
rect 76 644 82 647
rect 63 638 66 644
rect 82 638 85 644
rect 100 643 146 646
rect 153 644 156 651
rect 191 644 194 647
rect 211 644 214 647
rect 71 631 74 634
rect 91 631 94 634
rect 100 631 103 643
rect 153 641 184 644
rect 153 640 156 641
rect 191 641 214 644
rect 211 640 214 641
rect 124 632 127 636
rect 159 633 204 636
rect 211 636 212 640
rect 56 628 64 631
rect 71 628 103 631
rect 113 628 124 631
rect 39 596 43 599
rect 56 621 84 624
rect 56 599 59 621
rect 91 617 94 628
rect 62 605 65 613
rect 100 606 103 628
rect 120 618 124 621
rect 128 618 144 621
rect 125 612 128 618
rect 144 612 147 618
rect 133 605 136 608
rect 153 605 156 608
rect 159 605 162 633
rect 211 630 214 636
rect 104 602 126 605
rect 133 602 162 605
rect 5 549 8 596
rect 43 583 46 596
rect 58 598 59 599
rect 58 595 146 598
rect 153 591 156 602
rect 124 583 127 587
rect 182 583 185 626
rect 195 612 206 613
rect 220 615 223 667
rect 305 661 308 667
rect 324 661 327 667
rect 363 661 366 667
rect 366 657 382 660
rect 313 654 316 657
rect 333 654 336 657
rect 239 651 306 654
rect 236 631 239 651
rect 313 651 336 654
rect 363 651 366 657
rect 382 651 385 657
rect 246 644 252 647
rect 256 644 262 647
rect 243 638 246 644
rect 262 638 265 644
rect 280 643 326 646
rect 333 644 336 651
rect 371 644 374 647
rect 391 644 394 647
rect 251 631 254 634
rect 271 631 274 634
rect 280 631 283 643
rect 333 641 364 644
rect 333 640 336 641
rect 371 641 394 644
rect 391 640 394 641
rect 304 632 307 636
rect 339 633 384 636
rect 391 636 392 640
rect 236 628 244 631
rect 251 628 283 631
rect 293 628 304 631
rect 210 612 223 615
rect 236 621 264 624
rect 236 613 239 621
rect 271 617 274 628
rect 195 610 209 612
rect 195 606 198 610
rect 238 608 239 613
rect 207 602 209 606
rect 192 594 198 597
rect 206 597 209 602
rect 236 598 239 608
rect 242 605 245 613
rect 280 606 283 628
rect 300 618 304 621
rect 308 618 324 621
rect 305 612 308 618
rect 324 612 327 618
rect 313 605 316 608
rect 333 605 336 608
rect 339 605 342 633
rect 391 630 394 636
rect 284 602 306 605
rect 313 602 342 605
rect 206 593 207 597
rect 236 595 326 598
rect 206 590 209 593
rect 333 591 336 602
rect 208 586 209 590
rect 194 583 197 586
rect 304 583 307 587
rect 362 583 365 626
rect 399 623 402 667
rect 432 669 605 672
rect 609 669 649 672
rect 653 669 657 672
rect 661 669 677 672
rect 681 669 715 672
rect 719 669 785 672
rect 789 669 829 672
rect 833 669 837 672
rect 841 669 857 672
rect 861 669 895 672
rect 899 669 934 672
rect 432 623 435 669
rect 658 663 661 669
rect 677 663 680 669
rect 716 663 719 669
rect 719 659 735 662
rect 589 653 639 656
rect 666 656 669 659
rect 686 656 689 659
rect 643 653 659 656
rect 589 633 592 653
rect 666 653 689 656
rect 716 653 719 659
rect 735 653 738 659
rect 599 646 605 649
rect 609 646 615 649
rect 596 640 599 646
rect 615 640 618 646
rect 633 645 679 648
rect 686 646 689 653
rect 724 646 727 649
rect 744 646 747 649
rect 604 633 607 636
rect 624 633 627 636
rect 633 633 636 645
rect 686 643 717 646
rect 686 642 689 643
rect 724 643 747 646
rect 744 642 747 643
rect 657 634 660 638
rect 692 635 737 638
rect 744 638 745 642
rect 589 630 597 633
rect 604 630 636 633
rect 646 630 657 633
rect 589 623 617 626
rect 399 620 405 623
rect 375 612 386 613
rect 399 615 402 620
rect 390 612 402 615
rect 409 620 440 623
rect 405 614 408 619
rect 440 614 443 619
rect 375 610 389 612
rect 375 606 378 610
rect 387 605 389 606
rect 387 602 423 605
rect 372 594 378 597
rect 386 590 389 602
rect 399 593 407 596
rect 430 596 433 610
rect 414 593 444 596
rect 451 596 454 610
rect 589 601 592 623
rect 624 619 627 630
rect 595 607 598 615
rect 633 608 636 630
rect 653 620 657 623
rect 661 620 677 623
rect 658 614 661 620
rect 677 614 680 620
rect 666 607 669 610
rect 686 607 689 610
rect 692 607 695 635
rect 744 632 747 638
rect 637 604 659 607
rect 666 604 695 607
rect 591 600 592 601
rect 591 597 679 600
rect 451 593 464 596
rect 686 593 689 604
rect 414 590 417 593
rect 430 590 433 593
rect 451 590 454 593
rect 388 586 389 590
rect 374 583 377 586
rect 405 583 408 586
rect 421 583 424 586
rect 441 583 444 586
rect 66 580 84 583
rect 88 580 110 583
rect 114 580 124 583
rect 128 580 152 583
rect 156 580 181 583
rect 185 582 242 583
rect 185 580 204 582
rect 31 557 34 563
rect 18 554 35 557
rect 8 545 14 548
rect 5 533 8 545
rect 21 541 24 547
rect 43 548 46 579
rect 208 580 242 582
rect 246 580 264 583
rect 268 580 290 583
rect 294 580 304 583
rect 308 580 332 583
rect 336 580 361 583
rect 365 582 444 583
rect 365 580 384 582
rect 388 580 417 582
rect 421 580 444 582
rect 222 568 395 571
rect 434 561 437 580
rect 461 571 464 593
rect 657 585 660 589
rect 715 585 718 628
rect 728 614 739 615
rect 753 617 756 669
rect 838 663 841 669
rect 857 663 860 669
rect 896 663 899 669
rect 899 659 915 662
rect 769 654 816 656
rect 846 656 849 659
rect 866 656 869 659
rect 820 654 839 656
rect 769 653 839 654
rect 769 633 772 653
rect 846 653 869 656
rect 896 653 899 659
rect 915 653 918 659
rect 779 646 785 649
rect 789 646 795 649
rect 776 640 779 646
rect 795 640 798 646
rect 813 645 859 648
rect 866 646 869 653
rect 904 646 907 649
rect 924 646 927 649
rect 784 633 787 636
rect 804 633 807 636
rect 813 633 816 645
rect 866 643 897 646
rect 866 642 869 643
rect 904 643 927 646
rect 837 634 840 638
rect 872 635 917 638
rect 769 630 777 633
rect 784 630 816 633
rect 826 630 837 633
rect 743 614 756 617
rect 769 623 797 626
rect 769 615 772 623
rect 804 619 807 630
rect 728 612 742 614
rect 728 608 731 612
rect 771 610 772 615
rect 740 604 742 608
rect 725 596 731 599
rect 739 599 742 604
rect 769 600 772 610
rect 775 607 778 615
rect 813 608 816 630
rect 833 620 837 623
rect 841 620 857 623
rect 838 614 841 620
rect 857 614 860 620
rect 846 607 849 610
rect 866 607 869 610
rect 872 607 875 635
rect 924 632 927 643
rect 817 604 839 607
rect 846 604 875 607
rect 739 595 740 599
rect 769 597 859 600
rect 739 592 742 595
rect 866 593 869 604
rect 741 588 742 592
rect 727 585 730 588
rect 837 585 840 589
rect 895 585 898 628
rect 931 625 934 669
rect 931 622 937 625
rect 908 614 919 615
rect 931 617 934 622
rect 923 614 934 617
rect 941 622 972 625
rect 937 616 940 621
rect 972 616 975 621
rect 908 612 922 614
rect 908 608 911 612
rect 920 607 922 608
rect 920 604 955 607
rect 905 596 911 599
rect 919 592 922 604
rect 932 595 939 598
rect 962 598 965 612
rect 946 595 976 598
rect 946 592 949 595
rect 962 592 965 595
rect 983 592 986 612
rect 921 588 922 592
rect 907 585 910 588
rect 937 585 940 588
rect 953 585 956 588
rect 973 585 976 588
rect 599 582 617 585
rect 621 582 643 585
rect 647 582 657 585
rect 661 582 685 585
rect 689 582 714 585
rect 718 584 775 585
rect 718 582 737 584
rect 595 561 598 581
rect 741 582 775 584
rect 779 582 797 585
rect 801 582 823 585
rect 827 582 837 585
rect 841 582 865 585
rect 869 582 894 585
rect 898 584 976 585
rect 898 582 917 584
rect 921 582 949 584
rect 953 582 976 584
rect 755 570 928 573
rect 434 558 598 561
rect 39 545 43 548
rect 18 538 35 541
rect 8 529 14 532
rect 5 513 8 529
rect 21 521 24 538
rect 18 518 24 521
rect 8 510 14 513
rect 44 513 47 544
rect 983 536 986 588
rect 722 533 986 536
rect 39 509 43 512
rect 267 512 307 515
rect 311 512 315 515
rect 319 512 335 515
rect 339 512 373 515
rect 377 512 443 515
rect 447 512 487 515
rect 491 512 495 515
rect 499 512 515 515
rect 519 512 553 515
rect 557 512 592 515
rect 5 461 8 509
rect 31 469 34 474
rect 19 466 36 469
rect 9 457 15 460
rect 6 445 9 457
rect 22 453 25 459
rect 44 460 47 509
rect 316 506 319 512
rect 335 506 338 512
rect 374 506 377 512
rect 377 502 393 505
rect 324 499 327 502
rect 344 499 347 502
rect 250 496 317 499
rect 247 476 250 496
rect 324 496 347 499
rect 374 496 377 502
rect 393 496 396 502
rect 257 489 263 492
rect 267 489 273 492
rect 254 483 257 489
rect 273 483 276 489
rect 291 488 337 491
rect 344 489 347 496
rect 382 489 385 492
rect 402 489 405 492
rect 262 476 265 479
rect 282 476 285 479
rect 291 476 294 488
rect 344 486 375 489
rect 344 485 347 486
rect 382 486 405 489
rect 402 485 405 486
rect 315 477 318 481
rect 350 478 395 481
rect 402 481 403 485
rect 247 473 255 476
rect 262 473 294 476
rect 304 473 315 476
rect 247 466 275 469
rect 40 457 44 460
rect 19 450 36 453
rect 9 441 15 444
rect 6 425 9 441
rect 22 433 25 450
rect 19 430 25 433
rect 45 428 48 456
rect 247 443 250 466
rect 282 462 285 473
rect 253 450 256 458
rect 291 451 294 473
rect 311 463 315 466
rect 319 463 335 466
rect 316 457 319 463
rect 335 457 338 463
rect 324 450 327 453
rect 344 450 347 453
rect 350 450 353 478
rect 402 475 405 481
rect 295 447 317 450
rect 324 447 353 450
rect 249 440 337 443
rect 344 436 347 447
rect 315 428 318 432
rect 373 428 376 471
rect 386 457 397 458
rect 411 460 414 512
rect 496 506 499 512
rect 515 506 518 512
rect 554 506 557 512
rect 557 502 573 505
rect 504 499 507 502
rect 524 499 527 502
rect 431 496 497 499
rect 427 476 430 496
rect 504 496 527 499
rect 554 496 557 502
rect 573 496 576 502
rect 437 489 443 492
rect 447 489 453 492
rect 434 483 437 489
rect 453 483 456 489
rect 471 488 517 491
rect 524 489 527 496
rect 562 489 565 492
rect 582 489 585 492
rect 442 476 445 479
rect 462 476 465 479
rect 471 476 474 488
rect 524 486 555 489
rect 524 485 527 486
rect 562 486 585 489
rect 582 485 585 486
rect 495 477 498 481
rect 530 478 575 481
rect 427 473 435 476
rect 442 473 474 476
rect 484 473 495 476
rect 401 457 414 460
rect 427 466 455 469
rect 427 458 430 466
rect 462 462 465 473
rect 386 455 400 457
rect 386 451 389 455
rect 429 453 430 458
rect 398 447 400 451
rect 383 439 389 442
rect 397 442 400 447
rect 427 443 430 453
rect 433 450 436 458
rect 471 451 474 473
rect 491 463 495 466
rect 499 463 515 466
rect 496 457 499 463
rect 515 457 518 463
rect 504 450 507 453
rect 524 450 527 453
rect 530 450 533 478
rect 582 475 585 481
rect 475 447 497 450
rect 504 447 533 450
rect 397 438 398 442
rect 427 440 517 443
rect 397 435 400 438
rect 524 436 527 447
rect 399 431 400 435
rect 385 428 388 431
rect 495 428 498 432
rect 553 428 556 471
rect 589 468 592 512
rect 589 465 595 468
rect 566 457 577 458
rect 589 460 592 465
rect 581 457 592 460
rect 599 465 630 468
rect 595 459 598 464
rect 630 459 633 464
rect 566 455 580 457
rect 566 451 569 455
rect 578 450 580 451
rect 578 447 613 450
rect 563 439 569 442
rect 577 435 580 447
rect 590 438 597 441
rect 620 441 623 455
rect 604 438 634 441
rect 604 435 607 438
rect 620 435 623 438
rect 641 435 644 455
rect 579 431 580 435
rect 565 428 568 431
rect 595 428 598 431
rect 611 428 614 431
rect 631 428 634 431
rect 9 422 15 425
rect 44 425 253 428
rect 40 421 44 424
rect 257 425 275 428
rect 279 425 301 428
rect 305 425 315 428
rect 319 425 343 428
rect 347 425 372 428
rect 376 427 433 428
rect 376 425 395 427
rect 399 425 433 427
rect 437 425 455 428
rect 459 425 481 428
rect 485 425 495 428
rect 499 425 523 428
rect 527 425 552 428
rect 556 427 634 428
rect 556 425 575 427
rect 579 425 607 427
rect 611 425 634 427
rect 6 415 9 421
rect 6 380 9 411
rect 32 388 35 394
rect 20 385 37 388
rect 10 376 16 379
rect 7 364 10 376
rect 23 372 26 378
rect 45 379 48 421
rect 97 411 137 414
rect 141 411 145 414
rect 149 411 165 414
rect 169 411 203 414
rect 207 411 242 414
rect 413 413 586 416
rect 146 405 149 411
rect 165 405 168 411
rect 204 405 207 411
rect 207 401 223 404
rect 154 398 157 401
rect 174 398 177 401
rect 77 397 147 398
rect 62 395 147 397
rect 62 394 80 395
rect 154 395 177 398
rect 204 395 207 401
rect 223 395 226 401
rect 41 376 45 379
rect 20 369 37 372
rect 10 360 16 363
rect 7 344 10 360
rect 23 352 26 369
rect 20 349 26 352
rect 10 341 16 344
rect 46 344 49 375
rect 77 375 80 394
rect 87 388 93 391
rect 97 388 103 391
rect 84 382 87 388
rect 103 382 106 388
rect 121 387 167 390
rect 174 388 177 395
rect 212 388 215 391
rect 232 388 235 391
rect 92 375 95 378
rect 112 375 115 378
rect 121 375 124 387
rect 174 385 205 388
rect 174 384 177 385
rect 212 386 235 388
rect 212 385 232 386
rect 145 376 148 380
rect 180 377 225 380
rect 77 372 85 375
rect 92 372 124 375
rect 134 372 145 375
rect 41 340 45 343
rect 7 296 10 340
rect 46 327 49 340
rect 77 365 105 368
rect 77 342 80 365
rect 112 361 115 372
rect 83 349 86 357
rect 121 350 124 372
rect 141 362 145 365
rect 149 362 165 365
rect 146 356 149 362
rect 165 356 168 362
rect 154 349 157 352
rect 174 349 177 352
rect 180 349 183 377
rect 232 374 235 382
rect 125 346 147 349
rect 154 346 183 349
rect 239 380 242 411
rect 641 406 644 431
rect 722 394 725 533
rect 239 377 510 380
rect 514 377 554 380
rect 558 377 562 380
rect 566 377 582 380
rect 586 377 620 380
rect 624 377 690 380
rect 694 377 734 380
rect 738 377 742 380
rect 746 377 762 380
rect 766 377 800 380
rect 804 377 839 380
rect 77 339 167 342
rect 32 304 35 309
rect 20 301 37 304
rect 10 292 16 295
rect 7 280 10 292
rect 23 288 26 294
rect 46 295 49 323
rect 77 314 80 339
rect 174 335 177 346
rect 145 327 148 331
rect 203 327 206 370
rect 216 356 227 357
rect 239 359 242 377
rect 563 371 566 377
rect 582 371 585 377
rect 621 371 624 377
rect 624 367 640 370
rect 231 356 242 359
rect 494 361 541 364
rect 571 364 574 367
rect 591 364 594 367
rect 545 361 564 364
rect 216 354 230 356
rect 216 350 219 354
rect 228 346 230 350
rect 213 338 219 341
rect 227 340 230 346
rect 227 337 273 340
rect 227 334 230 337
rect 494 341 497 361
rect 571 361 594 364
rect 621 361 624 367
rect 640 361 643 367
rect 504 354 510 357
rect 514 354 520 357
rect 501 348 504 354
rect 520 348 523 354
rect 538 353 584 356
rect 591 354 594 361
rect 629 354 632 357
rect 649 354 652 357
rect 509 341 512 344
rect 529 341 532 344
rect 538 341 541 353
rect 591 351 622 354
rect 591 350 594 351
rect 629 351 652 354
rect 649 350 652 351
rect 562 342 565 346
rect 597 343 642 346
rect 649 346 650 350
rect 494 338 502 341
rect 509 338 541 341
rect 551 338 562 341
rect 229 330 230 334
rect 494 331 522 334
rect 215 327 218 330
rect 87 324 105 327
rect 109 324 131 327
rect 135 324 145 327
rect 149 324 173 327
rect 177 324 202 327
rect 206 326 453 327
rect 206 324 225 326
rect 229 324 453 326
rect 41 292 45 295
rect 20 285 37 288
rect 10 276 16 279
rect 7 260 10 276
rect 23 268 26 285
rect 20 265 26 268
rect 10 257 16 260
rect 46 260 49 291
rect 450 293 453 324
rect 494 309 497 331
rect 529 327 532 338
rect 500 315 503 323
rect 538 316 541 338
rect 558 328 562 331
rect 566 328 582 331
rect 563 322 566 328
rect 582 322 585 328
rect 571 315 574 318
rect 591 315 594 318
rect 597 315 600 343
rect 649 340 652 346
rect 542 312 564 315
rect 571 312 600 315
rect 478 308 497 309
rect 478 305 584 308
rect 591 301 594 312
rect 562 293 565 297
rect 620 293 623 336
rect 633 322 644 323
rect 658 325 661 377
rect 743 371 746 377
rect 762 371 765 377
rect 801 371 804 377
rect 804 367 820 370
rect 674 361 721 364
rect 751 364 754 367
rect 771 364 774 367
rect 725 361 744 364
rect 674 341 677 361
rect 751 361 774 364
rect 801 361 804 367
rect 820 361 823 367
rect 684 354 690 357
rect 694 354 700 357
rect 681 348 684 354
rect 700 348 703 354
rect 718 353 764 356
rect 771 354 774 361
rect 809 354 812 357
rect 829 354 832 357
rect 689 341 692 344
rect 709 341 712 344
rect 718 341 721 353
rect 771 351 802 354
rect 771 350 774 351
rect 809 351 832 354
rect 742 342 745 346
rect 777 343 822 346
rect 674 338 682 341
rect 689 338 721 341
rect 731 338 742 341
rect 648 322 661 325
rect 674 331 702 334
rect 674 323 677 331
rect 709 327 712 338
rect 633 320 647 322
rect 633 316 636 320
rect 676 318 677 323
rect 645 312 647 316
rect 630 304 636 307
rect 644 307 647 312
rect 674 308 677 318
rect 680 315 683 323
rect 718 316 721 338
rect 738 328 742 331
rect 746 328 762 331
rect 743 322 746 328
rect 762 322 765 328
rect 751 315 754 318
rect 771 315 774 318
rect 777 315 780 343
rect 829 340 832 351
rect 722 312 744 315
rect 751 312 780 315
rect 644 303 645 307
rect 674 305 764 308
rect 644 300 647 303
rect 771 301 774 312
rect 646 296 647 300
rect 632 293 635 296
rect 742 293 745 297
rect 800 293 803 336
rect 836 333 839 377
rect 836 330 842 333
rect 813 322 824 323
rect 836 325 839 330
rect 828 322 839 325
rect 846 330 877 333
rect 842 324 845 329
rect 877 324 880 329
rect 813 320 827 322
rect 813 316 816 320
rect 825 315 827 316
rect 825 312 860 315
rect 810 304 816 307
rect 824 300 827 312
rect 837 303 844 306
rect 867 306 870 320
rect 851 303 881 306
rect 851 300 854 303
rect 867 300 870 303
rect 888 300 891 320
rect 826 296 827 300
rect 812 293 815 296
rect 842 293 845 296
rect 858 293 861 296
rect 878 293 881 296
rect 450 290 500 293
rect 504 290 522 293
rect 526 290 548 293
rect 552 290 562 293
rect 566 290 590 293
rect 594 290 619 293
rect 623 292 680 293
rect 623 290 642 292
rect 646 290 680 292
rect 684 290 702 293
rect 706 290 728 293
rect 732 290 742 293
rect 746 290 770 293
rect 774 290 799 293
rect 803 292 881 293
rect 803 290 822 292
rect 826 290 854 292
rect 858 290 881 292
rect 660 278 833 281
rect 41 256 45 259
rect 888 259 891 296
rect 702 256 891 259
rect 7 238 10 256
rect 7 209 10 234
rect 32 217 35 223
rect 20 214 37 217
rect 10 205 16 208
rect 7 193 10 205
rect 23 201 26 207
rect 45 208 48 256
rect 114 225 154 228
rect 158 225 162 228
rect 166 225 182 228
rect 186 225 220 228
rect 224 225 290 228
rect 294 225 334 228
rect 338 225 342 228
rect 346 225 362 228
rect 366 225 400 228
rect 404 225 439 228
rect 74 212 77 224
rect 163 219 166 225
rect 182 219 185 225
rect 221 219 224 225
rect 224 215 240 218
rect 171 212 174 215
rect 191 212 194 215
rect 74 209 164 212
rect 41 205 45 208
rect 20 198 37 201
rect 10 189 16 192
rect 7 173 10 189
rect 23 181 26 198
rect 20 178 26 181
rect 10 170 16 173
rect 46 173 49 204
rect 94 189 97 209
rect 171 209 194 212
rect 221 209 224 215
rect 240 209 243 215
rect 104 202 110 205
rect 114 202 120 205
rect 101 196 104 202
rect 120 196 123 202
rect 138 201 184 204
rect 191 202 194 209
rect 229 202 232 205
rect 249 202 252 205
rect 109 189 112 192
rect 129 189 132 192
rect 138 189 141 201
rect 191 199 222 202
rect 191 198 194 199
rect 229 199 252 202
rect 249 198 252 199
rect 162 190 165 194
rect 197 191 242 194
rect 249 194 250 198
rect 94 186 102 189
rect 109 186 141 189
rect 151 186 162 189
rect 41 169 45 172
rect 7 121 10 169
rect 33 129 36 135
rect 46 129 49 169
rect 94 179 122 182
rect 94 156 97 179
rect 129 175 132 186
rect 100 163 103 171
rect 138 164 141 186
rect 158 176 162 179
rect 166 176 182 179
rect 163 170 166 176
rect 182 170 185 176
rect 171 163 174 166
rect 191 163 194 166
rect 197 163 200 191
rect 249 188 252 194
rect 142 160 164 163
rect 171 160 200 163
rect 74 153 184 156
rect 74 140 77 153
rect 191 149 194 160
rect 162 141 165 145
rect 220 141 223 184
rect 233 170 244 171
rect 258 173 261 225
rect 343 219 346 225
rect 362 219 365 225
rect 401 219 404 225
rect 404 215 420 218
rect 351 212 354 215
rect 371 212 374 215
rect 277 209 344 212
rect 274 189 277 209
rect 351 209 374 212
rect 401 209 404 215
rect 420 209 423 215
rect 284 202 290 205
rect 294 202 300 205
rect 281 196 284 202
rect 300 196 303 202
rect 318 201 364 204
rect 371 202 374 209
rect 409 202 412 205
rect 429 202 432 205
rect 289 189 292 192
rect 309 189 312 192
rect 318 189 321 201
rect 371 199 402 202
rect 371 198 374 199
rect 409 201 432 202
rect 409 199 429 201
rect 342 190 345 194
rect 377 191 422 194
rect 274 186 282 189
rect 289 186 321 189
rect 331 186 342 189
rect 248 170 261 173
rect 274 179 302 182
rect 274 171 277 179
rect 309 175 312 186
rect 233 168 247 170
rect 233 164 236 168
rect 276 166 277 171
rect 245 160 247 164
rect 230 152 236 155
rect 244 155 247 160
rect 274 156 277 166
rect 280 163 283 171
rect 318 164 321 186
rect 338 176 342 179
rect 346 176 362 179
rect 343 170 346 176
rect 362 170 365 176
rect 351 163 354 166
rect 371 163 374 166
rect 377 163 380 191
rect 429 188 432 197
rect 322 160 344 163
rect 351 160 380 163
rect 244 151 245 155
rect 274 153 364 156
rect 244 148 247 151
rect 371 149 374 160
rect 246 144 247 148
rect 232 141 235 144
rect 342 141 345 145
rect 400 141 403 184
rect 436 181 439 225
rect 436 178 442 181
rect 413 170 424 171
rect 436 173 439 178
rect 428 170 439 173
rect 446 178 477 181
rect 481 178 533 181
rect 537 178 577 181
rect 581 178 585 181
rect 589 178 605 181
rect 609 178 643 181
rect 647 178 713 181
rect 717 178 757 181
rect 761 178 765 181
rect 769 178 785 181
rect 789 178 823 181
rect 827 178 862 181
rect 442 172 445 177
rect 477 172 480 177
rect 586 172 589 178
rect 605 172 608 178
rect 644 172 647 178
rect 413 168 427 170
rect 647 168 663 171
rect 413 164 416 168
rect 425 163 427 164
rect 425 160 460 163
rect 410 152 416 155
rect 424 148 427 160
rect 437 151 444 154
rect 467 154 470 168
rect 488 165 491 168
rect 594 165 597 168
rect 614 165 617 168
rect 488 162 587 165
rect 451 151 481 154
rect 451 148 454 151
rect 467 148 470 151
rect 488 148 491 162
rect 426 144 427 148
rect 412 141 415 144
rect 442 141 445 144
rect 458 141 461 144
rect 478 141 481 144
rect 517 142 520 162
rect 594 162 617 165
rect 644 162 647 168
rect 663 162 666 168
rect 527 155 533 158
rect 537 155 543 158
rect 524 149 527 155
rect 543 149 546 155
rect 561 154 607 157
rect 614 155 617 162
rect 652 155 655 158
rect 672 155 675 158
rect 532 142 535 145
rect 552 142 555 145
rect 561 142 564 154
rect 614 152 645 155
rect 614 151 617 152
rect 652 152 675 155
rect 672 151 675 152
rect 585 143 588 147
rect 620 144 665 147
rect 672 147 673 151
rect 104 138 122 141
rect 126 138 148 141
rect 152 138 162 141
rect 166 138 190 141
rect 194 138 219 141
rect 223 140 280 141
rect 223 138 242 140
rect 100 129 103 137
rect 246 138 280 140
rect 284 138 302 141
rect 306 138 328 141
rect 332 138 342 141
rect 346 138 370 141
rect 374 138 399 141
rect 403 140 495 141
rect 403 138 422 140
rect 426 138 454 140
rect 458 138 495 140
rect 517 139 525 142
rect 532 139 564 142
rect 574 139 585 142
rect 21 126 38 129
rect 46 126 103 129
rect 260 126 433 129
rect 11 117 17 120
rect 8 105 11 117
rect 24 113 27 119
rect 46 120 49 126
rect 42 117 46 120
rect 21 110 38 113
rect 11 101 17 104
rect 8 85 11 101
rect 24 93 27 110
rect 21 90 27 93
rect 11 82 17 85
rect 47 85 50 116
rect 492 94 495 138
rect 517 132 545 135
rect 517 110 520 132
rect 552 128 555 139
rect 523 116 526 124
rect 561 117 564 139
rect 581 129 585 132
rect 589 129 605 132
rect 586 123 589 129
rect 605 123 608 129
rect 594 116 597 119
rect 614 116 617 119
rect 620 116 623 144
rect 672 141 675 147
rect 565 113 587 116
rect 594 113 623 116
rect 519 109 520 110
rect 519 106 607 109
rect 614 102 617 113
rect 585 94 588 98
rect 643 94 646 137
rect 656 123 667 124
rect 681 126 684 178
rect 766 172 769 178
rect 785 172 788 178
rect 824 172 827 178
rect 827 168 843 171
rect 774 165 777 168
rect 794 165 797 168
rect 701 162 767 165
rect 697 142 700 162
rect 774 162 797 165
rect 824 162 827 168
rect 843 162 846 168
rect 707 155 713 158
rect 717 155 723 158
rect 704 149 707 155
rect 723 149 726 155
rect 741 154 787 157
rect 794 155 797 162
rect 832 155 835 158
rect 852 155 855 158
rect 712 142 715 145
rect 732 142 735 145
rect 741 142 744 154
rect 794 152 825 155
rect 794 151 797 152
rect 832 152 855 155
rect 765 143 768 147
rect 800 144 845 147
rect 697 139 705 142
rect 712 139 744 142
rect 754 139 765 142
rect 671 123 684 126
rect 697 132 725 135
rect 697 124 700 132
rect 732 128 735 139
rect 656 121 670 123
rect 656 117 659 121
rect 699 119 700 124
rect 668 113 670 117
rect 653 105 659 108
rect 667 108 670 113
rect 697 109 700 119
rect 703 116 706 124
rect 741 117 744 139
rect 761 129 765 132
rect 769 129 785 132
rect 766 123 769 129
rect 785 123 788 129
rect 774 116 777 119
rect 794 116 797 119
rect 800 116 803 144
rect 852 141 855 152
rect 745 113 767 116
rect 774 113 803 116
rect 667 104 668 108
rect 697 106 787 109
rect 667 101 670 104
rect 794 102 797 113
rect 669 97 670 101
rect 655 94 658 97
rect 765 94 768 98
rect 823 94 826 137
rect 859 134 862 178
rect 859 131 865 134
rect 836 123 847 124
rect 859 126 862 131
rect 851 123 862 126
rect 869 131 900 134
rect 865 125 868 130
rect 900 125 903 130
rect 836 121 850 123
rect 836 117 839 121
rect 848 116 850 117
rect 848 113 883 116
rect 833 105 839 108
rect 847 101 850 113
rect 860 104 867 107
rect 890 107 893 121
rect 874 104 904 107
rect 874 101 877 104
rect 890 101 893 104
rect 911 101 914 121
rect 849 97 850 101
rect 835 94 838 97
rect 865 94 868 97
rect 881 94 884 97
rect 901 94 904 97
rect 492 91 523 94
rect 527 91 545 94
rect 549 91 571 94
rect 575 91 585 94
rect 589 91 613 94
rect 617 91 642 94
rect 646 93 703 94
rect 646 91 665 93
rect 669 91 703 93
rect 707 91 725 94
rect 729 91 751 94
rect 755 91 765 94
rect 769 91 793 94
rect 797 91 822 94
rect 826 93 904 94
rect 826 91 845 93
rect 849 91 877 93
rect 881 91 904 93
rect 42 81 46 84
rect 8 40 11 81
rect 33 48 36 54
rect 22 45 39 48
rect 12 36 18 39
rect 9 24 12 36
rect 25 32 28 38
rect 47 39 50 81
rect 683 79 856 82
rect 43 36 47 39
rect 22 29 39 32
rect 12 20 18 23
rect 9 4 12 20
rect 25 12 28 29
rect 22 9 28 12
rect 12 1 18 4
rect 48 4 51 35
rect 43 0 47 3
<< metal2 >>
rect 4 1259 87 1262
rect 30 1243 56 1246
rect 88 1240 91 1259
rect 77 1175 80 1193
rect 44 1172 77 1175
rect 116 1167 119 1194
rect 124 1175 127 1220
rect 132 1214 135 1259
rect 316 1241 319 1260
rect 124 1172 125 1175
rect 203 1167 206 1186
rect 116 1164 206 1167
rect 27 1158 70 1159
rect 31 1156 70 1158
rect 297 1088 301 1188
rect 305 1176 308 1194
rect 344 1168 347 1195
rect 352 1176 355 1221
rect 360 1215 363 1260
rect 352 1173 353 1176
rect 431 1168 434 1187
rect 456 1186 563 1189
rect 344 1165 434 1168
rect 297 1084 410 1088
rect 32 1073 241 1077
rect 6 1005 74 1008
rect 32 989 58 992
rect 75 986 78 1005
rect 56 906 59 933
rect 64 921 67 939
rect 103 913 106 940
rect 111 921 114 966
rect 119 960 122 1005
rect 238 993 241 1073
rect 255 986 258 1005
rect 218 974 233 977
rect 230 951 233 974
rect 230 948 235 951
rect 240 948 241 951
rect 111 918 112 921
rect 190 913 193 932
rect 213 932 223 935
rect 103 910 193 913
rect 220 910 223 932
rect 244 921 247 939
rect 283 913 286 940
rect 291 921 294 966
rect 299 960 302 1005
rect 407 980 410 1084
rect 560 991 563 1186
rect 570 983 573 1002
rect 398 977 410 980
rect 291 918 292 921
rect 370 913 373 932
rect 283 910 373 913
rect 398 910 401 931
rect 33 903 59 906
rect 441 900 469 904
rect 8 834 277 837
rect 33 815 264 818
rect 278 815 281 834
rect 35 734 239 737
rect 9 667 72 670
rect 35 651 55 654
rect 73 648 76 667
rect 55 583 58 595
rect 62 583 65 601
rect 47 580 62 583
rect 55 567 58 580
rect 101 575 104 602
rect 109 583 112 628
rect 117 622 120 667
rect 236 655 239 734
rect 260 721 263 762
rect 267 750 270 768
rect 306 742 309 769
rect 314 750 317 795
rect 322 789 325 834
rect 441 822 444 900
rect 552 895 555 930
rect 559 918 562 936
rect 598 910 601 937
rect 606 918 609 963
rect 614 957 617 1002
rect 606 915 607 918
rect 685 910 688 929
rect 598 907 688 910
rect 552 892 626 895
rect 458 815 461 834
rect 421 803 436 806
rect 433 780 436 803
rect 433 777 438 780
rect 443 777 444 780
rect 314 747 315 750
rect 393 742 396 761
rect 416 761 426 764
rect 306 739 396 742
rect 423 739 426 761
rect 447 750 450 768
rect 486 742 489 769
rect 494 750 497 795
rect 502 789 505 834
rect 623 810 626 892
rect 600 807 626 810
rect 494 747 495 750
rect 573 742 576 761
rect 486 739 576 742
rect 601 739 604 760
rect 260 717 410 721
rect 253 648 256 667
rect 216 636 231 639
rect 228 613 231 636
rect 228 610 233 613
rect 238 610 239 613
rect 109 580 110 583
rect 188 575 191 594
rect 211 594 221 597
rect 101 572 191 575
rect 218 572 221 594
rect 242 583 245 601
rect 281 575 284 602
rect 289 583 292 628
rect 297 622 300 667
rect 407 640 410 717
rect 606 650 609 669
rect 640 657 643 683
rect 396 637 410 640
rect 289 580 290 583
rect 368 575 371 594
rect 281 572 371 575
rect 396 572 399 593
rect 35 564 58 567
rect 427 566 460 569
rect 215 512 263 516
rect 215 506 218 512
rect 5 503 218 506
rect 231 496 246 499
rect 231 478 235 496
rect 264 493 267 512
rect 35 474 235 478
rect 10 411 93 414
rect 36 394 58 397
rect 94 392 97 411
rect 83 327 86 345
rect 50 323 83 326
rect 122 319 125 346
rect 130 327 133 372
rect 138 366 141 411
rect 246 386 249 439
rect 253 428 256 446
rect 292 420 295 447
rect 300 428 303 473
rect 308 467 311 512
rect 427 500 430 566
rect 587 552 590 597
rect 595 585 598 603
rect 634 577 637 604
rect 642 585 645 630
rect 650 624 653 669
rect 786 650 789 669
rect 817 658 820 691
rect 749 638 764 641
rect 761 615 764 638
rect 761 612 766 615
rect 771 612 772 615
rect 642 582 643 585
rect 721 577 724 596
rect 744 596 754 599
rect 634 574 724 577
rect 751 574 754 596
rect 775 585 778 603
rect 814 577 817 604
rect 822 585 825 630
rect 830 624 833 669
rect 822 582 823 585
rect 901 577 904 596
rect 814 574 904 577
rect 929 574 932 595
rect 587 549 618 552
rect 444 493 447 512
rect 407 481 422 484
rect 419 458 422 481
rect 419 455 424 458
rect 429 455 430 458
rect 300 425 301 428
rect 379 420 382 439
rect 402 439 412 442
rect 292 417 382 420
rect 409 417 412 439
rect 433 428 436 446
rect 472 420 475 447
rect 480 428 483 473
rect 488 467 491 512
rect 615 484 618 549
rect 586 481 618 484
rect 480 425 481 428
rect 559 420 562 439
rect 472 417 562 420
rect 587 417 590 438
rect 236 383 249 386
rect 542 402 640 405
rect 511 358 514 377
rect 542 365 545 402
rect 130 324 131 327
rect 209 319 212 338
rect 122 316 212 319
rect 36 310 76 312
rect 36 309 79 310
rect 10 234 113 237
rect 110 229 113 234
rect 36 224 73 227
rect 111 206 114 225
rect 100 141 103 159
rect 37 136 73 139
rect 139 133 142 160
rect 147 141 150 186
rect 155 180 158 225
rect 274 213 277 336
rect 291 206 294 225
rect 254 194 269 197
rect 266 171 269 194
rect 266 168 271 171
rect 276 168 277 171
rect 147 138 148 141
rect 226 133 229 152
rect 249 152 259 155
rect 139 130 229 133
rect 256 130 259 152
rect 280 141 283 159
rect 319 133 322 160
rect 327 141 330 186
rect 335 180 338 225
rect 472 201 476 305
rect 500 293 503 311
rect 539 285 542 312
rect 547 293 550 338
rect 555 332 558 377
rect 691 358 694 377
rect 722 365 725 390
rect 654 346 669 349
rect 666 323 669 346
rect 666 320 671 323
rect 676 320 677 323
rect 547 290 548 293
rect 626 285 629 304
rect 649 304 659 307
rect 539 282 629 285
rect 656 282 659 304
rect 680 293 683 311
rect 719 285 722 312
rect 727 293 730 338
rect 735 332 738 377
rect 727 290 728 293
rect 806 285 809 304
rect 719 282 809 285
rect 834 282 837 303
rect 433 198 476 201
rect 534 159 537 178
rect 327 138 328 141
rect 406 133 409 152
rect 319 130 409 133
rect 434 130 437 151
rect 516 58 519 106
rect 523 94 526 112
rect 562 86 565 113
rect 570 94 573 139
rect 578 133 581 178
rect 697 166 700 256
rect 714 159 717 178
rect 677 147 692 150
rect 689 124 692 147
rect 689 121 694 124
rect 699 121 700 124
rect 570 91 571 94
rect 649 86 652 105
rect 672 105 682 108
rect 562 83 652 86
rect 679 83 682 105
rect 703 94 706 112
rect 742 86 745 113
rect 750 94 753 139
rect 758 133 761 178
rect 750 91 751 94
rect 829 86 832 105
rect 742 83 832 86
rect 857 83 860 104
rect 37 55 519 58
<< ntransistor >>
rect 32 1317 35 1319
rect 32 1301 35 1303
rect 32 1281 35 1283
rect 32 1230 35 1232
rect 144 1228 146 1231
rect 164 1228 166 1231
rect 32 1214 35 1216
rect 372 1229 374 1232
rect 392 1229 394 1232
rect 202 1218 204 1221
rect 222 1218 224 1221
rect 82 1205 84 1208
rect 102 1205 104 1208
rect 430 1219 432 1222
rect 450 1219 452 1222
rect 310 1206 312 1209
rect 330 1206 332 1209
rect 32 1194 35 1196
rect 144 1179 146 1182
rect 164 1179 166 1182
rect 215 1179 217 1182
rect 372 1180 374 1183
rect 392 1180 394 1183
rect 443 1180 445 1183
rect 33 1142 36 1144
rect 33 1126 36 1128
rect 33 1106 36 1108
rect 34 1061 37 1063
rect 34 1045 37 1047
rect 34 1025 37 1027
rect 34 977 37 979
rect 131 974 133 977
rect 151 974 153 977
rect 34 961 37 963
rect 311 974 313 977
rect 331 974 333 977
rect 189 964 191 967
rect 209 964 211 967
rect 69 951 71 954
rect 89 951 91 954
rect 626 971 628 974
rect 646 971 648 974
rect 369 964 371 967
rect 389 964 391 967
rect 249 951 251 954
rect 269 951 271 954
rect 684 961 686 964
rect 704 961 706 964
rect 564 948 566 951
rect 584 948 586 951
rect 34 941 37 943
rect 131 925 133 928
rect 151 925 153 928
rect 202 925 204 928
rect 311 925 313 928
rect 331 925 333 928
rect 382 925 384 928
rect 412 924 414 927
rect 428 924 430 927
rect 448 924 450 928
rect 626 922 628 925
rect 646 922 648 925
rect 697 922 699 925
rect 34 890 37 892
rect 34 874 37 876
rect 34 854 37 856
rect 35 802 38 804
rect 334 803 336 806
rect 354 803 356 806
rect 35 786 38 788
rect 514 803 516 806
rect 534 803 536 806
rect 392 793 394 796
rect 412 793 414 796
rect 272 780 274 783
rect 292 780 294 783
rect 572 793 574 796
rect 592 793 594 796
rect 452 780 454 783
rect 472 780 474 783
rect 35 766 38 768
rect 334 754 336 757
rect 354 754 356 757
rect 405 754 407 757
rect 514 754 516 757
rect 534 754 536 757
rect 585 754 587 757
rect 614 753 616 756
rect 630 753 632 756
rect 650 753 652 757
rect 36 721 39 723
rect 36 705 39 707
rect 36 685 39 687
rect 36 637 39 639
rect 129 636 131 639
rect 149 636 151 639
rect 36 621 39 623
rect 309 636 311 639
rect 329 636 331 639
rect 187 626 189 629
rect 207 626 209 629
rect 67 613 69 616
rect 87 613 89 616
rect 662 638 664 641
rect 682 638 684 641
rect 367 626 369 629
rect 387 626 389 629
rect 247 613 249 616
rect 267 613 269 616
rect 842 638 844 641
rect 862 638 864 641
rect 720 628 722 631
rect 740 628 742 631
rect 600 615 602 618
rect 620 615 622 618
rect 900 628 902 631
rect 920 628 922 631
rect 780 615 782 618
rect 800 615 802 618
rect 36 601 39 603
rect 129 587 131 590
rect 149 587 151 590
rect 200 587 202 590
rect 309 587 311 590
rect 329 587 331 590
rect 380 587 382 590
rect 410 586 412 589
rect 426 586 428 589
rect 446 586 448 590
rect 662 589 664 592
rect 682 589 684 592
rect 733 589 735 592
rect 842 589 844 592
rect 862 589 864 592
rect 913 589 915 592
rect 942 588 944 591
rect 958 588 960 591
rect 978 588 980 592
rect 36 550 39 552
rect 36 534 39 536
rect 36 514 39 516
rect 320 481 322 484
rect 340 481 342 484
rect 37 462 40 464
rect 500 481 502 484
rect 520 481 522 484
rect 378 471 380 474
rect 398 471 400 474
rect 258 458 260 461
rect 278 458 280 461
rect 558 471 560 474
rect 578 471 580 474
rect 438 458 440 461
rect 458 458 460 461
rect 37 446 40 448
rect 320 432 322 435
rect 340 432 342 435
rect 391 432 393 435
rect 500 432 502 435
rect 520 432 522 435
rect 571 432 573 435
rect 600 431 602 434
rect 616 431 618 434
rect 636 431 638 435
rect 37 426 40 428
rect 38 381 41 383
rect 150 380 152 383
rect 170 380 172 383
rect 38 365 41 367
rect 208 370 210 373
rect 228 370 230 373
rect 88 357 90 360
rect 108 357 110 360
rect 38 345 41 347
rect 567 346 569 349
rect 587 346 589 349
rect 150 331 152 334
rect 170 331 172 334
rect 221 331 223 334
rect 747 346 749 349
rect 767 346 769 349
rect 625 336 627 339
rect 645 336 647 339
rect 505 323 507 326
rect 525 323 527 326
rect 805 336 807 339
rect 825 336 827 339
rect 685 323 687 326
rect 705 323 707 326
rect 38 297 41 299
rect 567 297 569 300
rect 587 297 589 300
rect 638 297 640 300
rect 747 297 749 300
rect 767 297 769 300
rect 818 297 820 300
rect 847 296 849 299
rect 863 296 865 299
rect 883 296 885 300
rect 38 281 41 283
rect 38 261 41 263
rect 38 210 41 212
rect 38 194 41 196
rect 167 194 169 197
rect 187 194 189 197
rect 38 174 41 176
rect 347 194 349 197
rect 367 194 369 197
rect 225 184 227 187
rect 245 184 247 187
rect 105 171 107 174
rect 125 171 127 174
rect 405 184 407 187
rect 425 184 427 187
rect 285 171 287 174
rect 305 171 307 174
rect 167 145 169 148
rect 187 145 189 148
rect 238 145 240 148
rect 347 145 349 148
rect 367 145 369 148
rect 418 145 420 148
rect 447 144 449 147
rect 463 144 465 147
rect 483 144 485 148
rect 590 147 592 150
rect 610 147 612 150
rect 770 147 772 150
rect 790 147 792 150
rect 648 137 650 140
rect 668 137 670 140
rect 528 124 530 127
rect 548 124 550 127
rect 39 122 42 124
rect 828 137 830 140
rect 848 137 850 140
rect 708 124 710 127
rect 728 124 730 127
rect 39 106 42 108
rect 590 98 592 101
rect 610 98 612 101
rect 661 98 663 101
rect 770 98 772 101
rect 790 98 792 101
rect 841 98 843 101
rect 870 97 872 100
rect 886 97 888 100
rect 906 97 908 101
rect 39 86 42 88
rect 40 41 43 43
rect 40 25 43 27
rect 40 5 43 7
<< ptransistor >>
rect 9 1317 15 1319
rect 9 1301 15 1303
rect 9 1281 15 1283
rect 144 1248 146 1254
rect 164 1248 166 1254
rect 372 1249 374 1255
rect 392 1249 394 1255
rect 9 1230 15 1232
rect 82 1225 84 1231
rect 102 1225 104 1231
rect 202 1238 204 1244
rect 222 1238 224 1244
rect 9 1214 15 1216
rect 310 1226 312 1232
rect 330 1226 332 1232
rect 430 1239 432 1245
rect 450 1239 452 1245
rect 144 1199 146 1205
rect 164 1199 166 1205
rect 372 1200 374 1206
rect 392 1200 394 1206
rect 9 1194 15 1196
rect 215 1193 217 1199
rect 443 1194 445 1200
rect 10 1142 16 1144
rect 10 1126 16 1128
rect 10 1106 16 1108
rect 11 1061 17 1063
rect 11 1045 17 1047
rect 11 1025 17 1027
rect 131 994 133 1000
rect 151 994 153 1000
rect 311 994 313 1000
rect 331 994 333 1000
rect 11 977 17 979
rect 69 971 71 977
rect 89 971 91 977
rect 189 984 191 990
rect 209 984 211 990
rect 11 961 17 963
rect 249 971 251 977
rect 269 971 271 977
rect 626 991 628 997
rect 646 991 648 997
rect 369 984 371 990
rect 389 984 391 990
rect 131 945 133 951
rect 151 945 153 951
rect 564 968 566 974
rect 584 968 586 974
rect 684 981 686 987
rect 704 981 706 987
rect 311 945 313 951
rect 331 945 333 951
rect 412 947 414 953
rect 428 947 430 953
rect 448 947 450 953
rect 11 941 17 943
rect 202 939 204 945
rect 382 939 384 945
rect 626 942 628 948
rect 646 942 648 948
rect 697 936 699 942
rect 11 890 17 892
rect 11 874 17 876
rect 11 854 17 856
rect 334 823 336 829
rect 354 823 356 829
rect 514 823 516 829
rect 534 823 536 829
rect 12 802 18 804
rect 272 800 274 806
rect 292 800 294 806
rect 392 813 394 819
rect 412 813 414 819
rect 12 786 18 788
rect 452 800 454 806
rect 472 800 474 806
rect 572 813 574 819
rect 592 813 594 819
rect 334 774 336 780
rect 354 774 356 780
rect 514 774 516 780
rect 534 774 536 780
rect 614 776 616 782
rect 630 776 632 782
rect 650 776 652 782
rect 12 766 18 768
rect 405 768 407 774
rect 585 768 587 774
rect 13 721 19 723
rect 13 705 19 707
rect 13 685 19 687
rect 129 656 131 662
rect 149 656 151 662
rect 309 656 311 662
rect 329 656 331 662
rect 662 658 664 664
rect 682 658 684 664
rect 842 658 844 664
rect 862 658 864 664
rect 13 637 19 639
rect 67 633 69 639
rect 87 633 89 639
rect 187 646 189 652
rect 207 646 209 652
rect 13 621 19 623
rect 247 633 249 639
rect 267 633 269 639
rect 367 646 369 652
rect 387 646 389 652
rect 129 607 131 613
rect 149 607 151 613
rect 600 635 602 641
rect 620 635 622 641
rect 720 648 722 654
rect 740 648 742 654
rect 309 607 311 613
rect 329 607 331 613
rect 780 635 782 641
rect 800 635 802 641
rect 900 648 902 654
rect 920 648 922 654
rect 410 609 412 615
rect 426 609 428 615
rect 446 609 448 615
rect 662 609 664 615
rect 682 609 684 615
rect 842 609 844 615
rect 862 609 864 615
rect 942 611 944 617
rect 958 611 960 617
rect 978 611 980 617
rect 13 601 19 603
rect 200 601 202 607
rect 380 601 382 607
rect 733 603 735 609
rect 913 603 915 609
rect 13 550 19 552
rect 13 534 19 536
rect 13 514 19 516
rect 320 501 322 507
rect 340 501 342 507
rect 500 501 502 507
rect 520 501 522 507
rect 258 478 260 484
rect 278 478 280 484
rect 378 491 380 497
rect 398 491 400 497
rect 14 462 20 464
rect 438 478 440 484
rect 458 478 460 484
rect 558 491 560 497
rect 578 491 580 497
rect 320 452 322 458
rect 340 452 342 458
rect 500 452 502 458
rect 520 452 522 458
rect 600 454 602 460
rect 616 454 618 460
rect 636 454 638 460
rect 14 446 20 448
rect 391 446 393 452
rect 571 446 573 452
rect 14 426 20 428
rect 150 400 152 406
rect 170 400 172 406
rect 15 381 21 383
rect 88 377 90 383
rect 108 377 110 383
rect 208 390 210 396
rect 228 390 230 396
rect 15 365 21 367
rect 567 366 569 372
rect 587 366 589 372
rect 747 366 749 372
rect 767 366 769 372
rect 150 351 152 357
rect 170 351 172 357
rect 15 345 21 347
rect 221 345 223 351
rect 505 343 507 349
rect 525 343 527 349
rect 625 356 627 362
rect 645 356 647 362
rect 685 343 687 349
rect 705 343 707 349
rect 805 356 807 362
rect 825 356 827 362
rect 567 317 569 323
rect 587 317 589 323
rect 747 317 749 323
rect 767 317 769 323
rect 847 319 849 325
rect 863 319 865 325
rect 883 319 885 325
rect 15 297 21 299
rect 638 311 640 317
rect 818 311 820 317
rect 15 281 21 283
rect 15 261 21 263
rect 167 214 169 220
rect 187 214 189 220
rect 347 214 349 220
rect 367 214 369 220
rect 15 210 21 212
rect 15 194 21 196
rect 105 191 107 197
rect 125 191 127 197
rect 225 204 227 210
rect 245 204 247 210
rect 15 174 21 176
rect 285 191 287 197
rect 305 191 307 197
rect 405 204 407 210
rect 425 204 427 210
rect 167 165 169 171
rect 187 165 189 171
rect 347 165 349 171
rect 367 165 369 171
rect 447 167 449 173
rect 463 167 465 173
rect 483 167 485 173
rect 590 167 592 173
rect 610 167 612 173
rect 770 167 772 173
rect 790 167 792 173
rect 238 159 240 165
rect 418 159 420 165
rect 528 144 530 150
rect 548 144 550 150
rect 648 157 650 163
rect 668 157 670 163
rect 708 144 710 150
rect 728 144 730 150
rect 828 157 830 163
rect 848 157 850 163
rect 16 122 22 124
rect 590 118 592 124
rect 610 118 612 124
rect 770 118 772 124
rect 790 118 792 124
rect 870 120 872 126
rect 886 120 888 126
rect 906 120 908 126
rect 16 106 22 108
rect 661 112 663 118
rect 841 112 843 118
rect 16 86 22 88
rect 17 41 23 43
rect 17 25 23 27
rect 17 5 23 7
<< polycontact >>
rect 17 1314 21 1318
rect 24 1298 28 1302
rect 17 1278 21 1282
rect 141 1242 145 1246
rect 17 1227 21 1231
rect 161 1235 165 1239
rect 369 1243 373 1247
rect 199 1232 203 1236
rect 79 1219 83 1223
rect 24 1211 28 1215
rect 219 1225 223 1229
rect 389 1236 393 1240
rect 427 1233 431 1237
rect 307 1220 311 1224
rect 99 1212 103 1216
rect 447 1226 451 1230
rect 327 1213 331 1217
rect 17 1191 21 1195
rect 141 1193 145 1197
rect 369 1194 373 1198
rect 161 1186 165 1190
rect 213 1186 217 1190
rect 389 1187 393 1191
rect 441 1187 445 1191
rect 18 1139 22 1143
rect 25 1123 29 1127
rect 18 1103 22 1107
rect 19 1058 23 1062
rect 26 1042 30 1046
rect 19 1022 23 1026
rect 128 988 132 992
rect 19 974 23 978
rect 148 981 152 985
rect 308 988 312 992
rect 186 978 190 982
rect 66 965 70 969
rect 26 958 30 962
rect 206 971 210 975
rect 328 981 332 985
rect 623 985 627 989
rect 366 978 370 982
rect 246 965 250 969
rect 86 958 90 962
rect 386 971 390 975
rect 643 978 647 982
rect 681 975 685 979
rect 561 962 565 966
rect 266 958 270 962
rect 701 968 705 972
rect 581 955 585 959
rect 19 938 23 942
rect 128 939 132 943
rect 308 939 312 943
rect 148 932 152 936
rect 200 932 204 936
rect 328 932 332 936
rect 380 932 384 936
rect 425 940 429 944
rect 409 931 413 935
rect 623 936 627 940
rect 446 931 450 935
rect 643 929 647 933
rect 695 929 699 933
rect 19 887 23 891
rect 26 871 30 875
rect 19 851 23 855
rect 331 817 335 821
rect 20 799 24 803
rect 351 810 355 814
rect 511 817 515 821
rect 389 807 393 811
rect 269 794 273 798
rect 27 783 31 787
rect 409 800 413 804
rect 531 810 535 814
rect 569 807 573 811
rect 449 794 453 798
rect 289 787 293 791
rect 589 800 593 804
rect 469 787 473 791
rect 331 768 335 772
rect 20 763 24 767
rect 511 768 515 772
rect 351 761 355 765
rect 403 761 407 765
rect 531 761 535 765
rect 583 761 587 765
rect 627 769 631 773
rect 611 760 615 764
rect 648 760 652 764
rect 21 718 25 722
rect 28 702 32 706
rect 21 682 25 686
rect 126 650 130 654
rect 21 634 25 638
rect 146 643 150 647
rect 306 650 310 654
rect 184 640 188 644
rect 64 627 68 631
rect 28 618 32 622
rect 204 633 208 637
rect 659 652 663 656
rect 326 643 330 647
rect 364 640 368 644
rect 244 627 248 631
rect 84 620 88 624
rect 384 633 388 637
rect 679 645 683 649
rect 839 652 843 656
rect 717 642 721 646
rect 597 629 601 633
rect 264 620 268 624
rect 737 635 741 639
rect 859 645 863 649
rect 897 642 901 646
rect 777 629 781 633
rect 617 622 621 626
rect 917 635 921 639
rect 797 622 801 626
rect 21 598 25 602
rect 126 601 130 605
rect 306 601 310 605
rect 146 594 150 598
rect 198 594 202 598
rect 326 594 330 598
rect 378 594 382 598
rect 423 602 427 606
rect 407 593 411 597
rect 659 603 663 607
rect 444 593 448 597
rect 839 603 843 607
rect 679 596 683 600
rect 731 596 735 600
rect 859 596 863 600
rect 911 596 915 600
rect 955 604 959 608
rect 939 595 943 599
rect 976 595 980 599
rect 21 547 25 551
rect 28 531 32 535
rect 21 511 25 515
rect 317 495 321 499
rect 337 488 341 492
rect 497 495 501 499
rect 375 485 379 489
rect 255 472 259 476
rect 22 459 26 463
rect 395 478 399 482
rect 517 488 521 492
rect 555 485 559 489
rect 435 472 439 476
rect 275 465 279 469
rect 575 478 579 482
rect 455 465 459 469
rect 29 443 33 447
rect 317 446 321 450
rect 497 446 501 450
rect 337 439 341 443
rect 389 439 393 443
rect 517 439 521 443
rect 569 439 573 443
rect 613 447 617 451
rect 597 438 601 442
rect 634 438 638 442
rect 22 423 26 427
rect 147 394 151 398
rect 23 378 27 382
rect 167 387 171 391
rect 205 384 209 388
rect 85 371 89 375
rect 30 362 34 366
rect 225 377 229 381
rect 105 364 109 368
rect 564 360 568 364
rect 23 342 27 346
rect 147 345 151 349
rect 584 353 588 357
rect 744 360 748 364
rect 622 350 626 354
rect 167 338 171 342
rect 219 338 223 342
rect 502 337 506 341
rect 642 343 646 347
rect 764 353 768 357
rect 802 350 806 354
rect 682 337 686 341
rect 522 330 526 334
rect 822 343 826 347
rect 702 330 706 334
rect 564 311 568 315
rect 23 294 27 298
rect 744 311 748 315
rect 584 304 588 308
rect 636 304 640 308
rect 764 304 768 308
rect 816 304 820 308
rect 860 312 864 316
rect 844 303 848 307
rect 881 303 885 307
rect 30 278 34 282
rect 23 258 27 262
rect 23 207 27 211
rect 164 208 168 212
rect 30 191 34 195
rect 184 201 188 205
rect 344 208 348 212
rect 222 198 226 202
rect 102 185 106 189
rect 23 171 27 175
rect 242 191 246 195
rect 364 201 368 205
rect 402 198 406 202
rect 282 185 286 189
rect 122 178 126 182
rect 422 191 426 195
rect 302 178 306 182
rect 164 159 168 163
rect 344 159 348 163
rect 184 152 188 156
rect 236 152 240 156
rect 364 152 368 156
rect 416 152 420 156
rect 460 160 464 164
rect 444 151 448 155
rect 587 161 591 165
rect 481 151 485 155
rect 607 154 611 158
rect 767 161 771 165
rect 645 151 649 155
rect 525 138 529 142
rect 665 144 669 148
rect 787 154 791 158
rect 825 151 829 155
rect 705 138 709 142
rect 545 131 549 135
rect 24 119 28 123
rect 845 144 849 148
rect 725 131 729 135
rect 587 112 591 116
rect 31 103 35 107
rect 767 112 771 116
rect 607 105 611 109
rect 659 105 663 109
rect 787 105 791 109
rect 839 105 843 109
rect 883 113 887 117
rect 867 104 871 108
rect 904 104 908 108
rect 24 83 28 87
rect 25 38 29 42
rect 32 22 36 26
rect 25 2 29 6
<< ndcontact >>
rect 31 1320 35 1324
rect 31 1312 35 1316
rect 31 1304 35 1308
rect 31 1276 35 1280
rect 31 1233 35 1237
rect 31 1225 35 1229
rect 139 1228 143 1232
rect 167 1228 171 1232
rect 31 1217 35 1221
rect 77 1205 81 1209
rect 197 1218 201 1222
rect 367 1229 371 1233
rect 395 1229 399 1233
rect 225 1218 229 1222
rect 105 1205 109 1209
rect 305 1206 309 1210
rect 425 1219 429 1223
rect 453 1219 457 1223
rect 333 1206 337 1210
rect 31 1189 35 1193
rect 139 1179 143 1183
rect 167 1179 171 1183
rect 209 1178 213 1182
rect 219 1178 223 1182
rect 367 1180 371 1184
rect 395 1180 399 1184
rect 437 1179 441 1183
rect 447 1179 451 1183
rect 32 1145 36 1149
rect 32 1137 36 1141
rect 32 1129 36 1133
rect 32 1101 36 1105
rect 33 1064 37 1068
rect 33 1056 37 1060
rect 33 1048 37 1052
rect 33 1020 37 1024
rect 33 980 37 984
rect 33 972 37 976
rect 126 974 130 978
rect 154 974 158 978
rect 33 964 37 968
rect 64 951 68 955
rect 184 964 188 968
rect 306 974 310 978
rect 334 974 338 978
rect 212 964 216 968
rect 92 951 96 955
rect 244 951 248 955
rect 364 964 368 968
rect 621 971 625 975
rect 649 971 653 975
rect 392 964 396 968
rect 272 951 276 955
rect 559 948 563 952
rect 679 961 683 965
rect 707 961 711 965
rect 587 948 591 952
rect 33 936 37 940
rect 126 925 130 929
rect 154 925 158 929
rect 196 924 200 928
rect 206 924 210 928
rect 306 925 310 929
rect 334 925 338 929
rect 376 924 380 928
rect 386 924 390 928
rect 407 924 411 928
rect 415 924 419 928
rect 423 924 427 928
rect 431 924 435 928
rect 442 924 446 928
rect 452 924 456 928
rect 621 922 625 926
rect 649 922 653 926
rect 691 921 695 925
rect 701 921 705 925
rect 33 893 37 897
rect 33 885 37 889
rect 33 877 37 881
rect 33 849 37 853
rect 34 805 38 809
rect 34 797 38 801
rect 329 803 333 807
rect 357 803 361 807
rect 34 789 38 793
rect 267 780 271 784
rect 387 793 391 797
rect 509 803 513 807
rect 537 803 541 807
rect 415 793 419 797
rect 295 780 299 784
rect 447 780 451 784
rect 567 793 571 797
rect 595 793 599 797
rect 475 780 479 784
rect 34 761 38 765
rect 329 754 333 758
rect 357 754 361 758
rect 399 753 403 757
rect 409 753 413 757
rect 509 754 513 758
rect 537 754 541 758
rect 579 753 583 757
rect 589 753 593 757
rect 609 753 613 757
rect 617 753 621 757
rect 625 753 629 757
rect 633 753 637 757
rect 644 753 648 757
rect 654 753 658 757
rect 35 724 39 728
rect 35 716 39 720
rect 35 708 39 712
rect 35 680 39 684
rect 35 640 39 644
rect 35 632 39 636
rect 124 636 128 640
rect 152 636 156 640
rect 35 624 39 628
rect 62 613 66 617
rect 182 626 186 630
rect 304 636 308 640
rect 332 636 336 640
rect 210 626 214 630
rect 90 613 94 617
rect 242 613 246 617
rect 362 626 366 630
rect 657 638 661 642
rect 685 638 689 642
rect 390 626 394 630
rect 270 613 274 617
rect 595 615 599 619
rect 715 628 719 632
rect 837 638 841 642
rect 865 638 869 642
rect 743 628 747 632
rect 623 615 627 619
rect 775 615 779 619
rect 895 628 899 632
rect 923 628 927 632
rect 803 615 807 619
rect 35 596 39 600
rect 124 587 128 591
rect 152 587 156 591
rect 194 586 198 590
rect 204 586 208 590
rect 304 587 308 591
rect 332 587 336 591
rect 374 586 378 590
rect 384 586 388 590
rect 405 586 409 590
rect 413 586 417 590
rect 421 586 425 590
rect 429 586 433 590
rect 440 586 444 590
rect 450 586 454 590
rect 657 589 661 593
rect 685 589 689 593
rect 727 588 731 592
rect 737 588 741 592
rect 837 589 841 593
rect 865 589 869 593
rect 907 588 911 592
rect 917 588 921 592
rect 937 588 941 592
rect 945 588 949 592
rect 953 588 957 592
rect 961 588 965 592
rect 972 588 976 592
rect 982 588 986 592
rect 35 553 39 557
rect 35 545 39 549
rect 35 537 39 541
rect 35 509 39 513
rect 315 481 319 485
rect 343 481 347 485
rect 36 465 40 469
rect 36 457 40 461
rect 253 458 257 462
rect 373 471 377 475
rect 495 481 499 485
rect 523 481 527 485
rect 401 471 405 475
rect 281 458 285 462
rect 36 449 40 453
rect 433 458 437 462
rect 553 471 557 475
rect 581 471 585 475
rect 461 458 465 462
rect 315 432 319 436
rect 343 432 347 436
rect 385 431 389 435
rect 395 431 399 435
rect 495 432 499 436
rect 523 432 527 436
rect 565 431 569 435
rect 575 431 579 435
rect 595 431 599 435
rect 603 431 607 435
rect 611 431 615 435
rect 619 431 623 435
rect 630 431 634 435
rect 640 431 644 435
rect 36 421 40 425
rect 37 384 41 388
rect 37 376 41 380
rect 145 380 149 384
rect 173 380 177 384
rect 37 368 41 372
rect 83 357 87 361
rect 203 370 207 374
rect 231 370 235 374
rect 111 357 115 361
rect 37 340 41 344
rect 145 331 149 335
rect 562 346 566 350
rect 590 346 594 350
rect 173 331 177 335
rect 215 330 219 334
rect 225 330 229 334
rect 500 323 504 327
rect 620 336 624 340
rect 742 346 746 350
rect 770 346 774 350
rect 648 336 652 340
rect 528 323 532 327
rect 680 323 684 327
rect 800 336 804 340
rect 828 336 832 340
rect 708 323 712 327
rect 37 300 41 304
rect 562 297 566 301
rect 590 297 594 301
rect 37 292 41 296
rect 632 296 636 300
rect 642 296 646 300
rect 742 297 746 301
rect 770 297 774 301
rect 812 296 816 300
rect 822 296 826 300
rect 842 296 846 300
rect 850 296 854 300
rect 858 296 862 300
rect 866 296 870 300
rect 877 296 881 300
rect 887 296 891 300
rect 37 284 41 288
rect 37 256 41 260
rect 37 213 41 217
rect 37 205 41 209
rect 37 197 41 201
rect 162 194 166 198
rect 190 194 194 198
rect 37 169 41 173
rect 100 171 104 175
rect 220 184 224 188
rect 342 194 346 198
rect 370 194 374 198
rect 248 184 252 188
rect 128 171 132 175
rect 280 171 284 175
rect 400 184 404 188
rect 428 184 432 188
rect 308 171 312 175
rect 162 145 166 149
rect 190 145 194 149
rect 232 144 236 148
rect 242 144 246 148
rect 342 145 346 149
rect 370 145 374 149
rect 412 144 416 148
rect 422 144 426 148
rect 442 144 446 148
rect 450 144 454 148
rect 458 144 462 148
rect 466 144 470 148
rect 477 144 481 148
rect 487 144 491 148
rect 585 147 589 151
rect 613 147 617 151
rect 38 125 42 129
rect 523 124 527 128
rect 643 137 647 141
rect 765 147 769 151
rect 793 147 797 151
rect 671 137 675 141
rect 551 124 555 128
rect 38 117 42 121
rect 703 124 707 128
rect 823 137 827 141
rect 851 137 855 141
rect 731 124 735 128
rect 38 109 42 113
rect 585 98 589 102
rect 613 98 617 102
rect 655 97 659 101
rect 665 97 669 101
rect 765 98 769 102
rect 793 98 797 102
rect 835 97 839 101
rect 845 97 849 101
rect 865 97 869 101
rect 873 97 877 101
rect 881 97 885 101
rect 889 97 893 101
rect 900 97 904 101
rect 910 97 914 101
rect 38 81 42 85
rect 39 44 43 48
rect 39 36 43 40
rect 39 28 43 32
rect 39 0 43 4
<< pdcontact >>
rect 10 1321 14 1325
rect 10 1312 14 1316
rect 10 1304 14 1308
rect 10 1296 14 1300
rect 10 1284 14 1288
rect 10 1276 14 1280
rect 139 1249 143 1253
rect 147 1249 151 1253
rect 159 1249 163 1253
rect 167 1249 171 1253
rect 367 1250 371 1254
rect 375 1250 379 1254
rect 387 1250 391 1254
rect 395 1250 399 1254
rect 10 1234 14 1238
rect 10 1225 14 1229
rect 77 1226 81 1230
rect 85 1226 89 1230
rect 97 1226 101 1230
rect 105 1226 109 1230
rect 197 1239 201 1243
rect 205 1239 209 1243
rect 217 1239 221 1243
rect 225 1239 229 1243
rect 10 1217 14 1221
rect 10 1209 14 1213
rect 10 1197 14 1201
rect 305 1227 309 1231
rect 313 1227 317 1231
rect 325 1227 329 1231
rect 333 1227 337 1231
rect 425 1240 429 1244
rect 433 1240 437 1244
rect 445 1240 449 1244
rect 453 1240 457 1244
rect 139 1200 143 1204
rect 147 1200 151 1204
rect 159 1200 163 1204
rect 167 1200 171 1204
rect 367 1201 371 1205
rect 375 1201 379 1205
rect 387 1201 391 1205
rect 395 1201 399 1205
rect 10 1189 14 1193
rect 210 1194 214 1198
rect 218 1194 222 1198
rect 438 1195 442 1199
rect 446 1195 450 1199
rect 11 1146 15 1150
rect 11 1137 15 1141
rect 11 1129 15 1133
rect 11 1121 15 1125
rect 11 1109 15 1113
rect 11 1101 15 1105
rect 12 1065 16 1069
rect 12 1056 16 1060
rect 12 1048 16 1052
rect 12 1040 16 1044
rect 12 1028 16 1032
rect 12 1020 16 1024
rect 126 995 130 999
rect 134 995 138 999
rect 146 995 150 999
rect 154 995 158 999
rect 306 995 310 999
rect 314 995 318 999
rect 326 995 330 999
rect 334 995 338 999
rect 12 981 16 985
rect 12 972 16 976
rect 64 972 68 976
rect 72 972 76 976
rect 84 972 88 976
rect 92 972 96 976
rect 184 985 188 989
rect 192 985 196 989
rect 204 985 208 989
rect 212 985 216 989
rect 12 964 16 968
rect 12 956 16 960
rect 12 944 16 948
rect 244 972 248 976
rect 252 972 256 976
rect 264 972 268 976
rect 272 972 276 976
rect 621 992 625 996
rect 629 992 633 996
rect 641 992 645 996
rect 649 992 653 996
rect 364 985 368 989
rect 372 985 376 989
rect 384 985 388 989
rect 392 985 396 989
rect 126 946 130 950
rect 134 946 138 950
rect 146 946 150 950
rect 559 969 563 973
rect 567 969 571 973
rect 579 969 583 973
rect 587 969 591 973
rect 679 982 683 986
rect 687 982 691 986
rect 699 982 703 986
rect 707 982 711 986
rect 154 946 158 950
rect 306 946 310 950
rect 314 946 318 950
rect 326 946 330 950
rect 334 946 338 950
rect 407 948 411 952
rect 431 948 435 952
rect 442 948 446 952
rect 452 948 456 952
rect 12 936 16 940
rect 197 940 201 944
rect 205 940 209 944
rect 377 940 381 944
rect 385 940 389 944
rect 621 943 625 947
rect 629 943 633 947
rect 641 943 645 947
rect 649 943 653 947
rect 692 937 696 941
rect 700 937 704 941
rect 12 894 16 898
rect 12 885 16 889
rect 12 877 16 881
rect 12 869 16 873
rect 12 857 16 861
rect 12 849 16 853
rect 329 824 333 828
rect 337 824 341 828
rect 349 824 353 828
rect 357 824 361 828
rect 509 824 513 828
rect 517 824 521 828
rect 529 824 533 828
rect 537 824 541 828
rect 13 806 17 810
rect 13 797 17 801
rect 267 801 271 805
rect 275 801 279 805
rect 287 801 291 805
rect 295 801 299 805
rect 387 814 391 818
rect 395 814 399 818
rect 407 814 411 818
rect 415 814 419 818
rect 13 789 17 793
rect 13 781 17 785
rect 13 769 17 773
rect 447 801 451 805
rect 455 801 459 805
rect 467 801 471 805
rect 475 801 479 805
rect 567 814 571 818
rect 575 814 579 818
rect 587 814 591 818
rect 595 814 599 818
rect 329 775 333 779
rect 337 775 341 779
rect 349 775 353 779
rect 357 775 361 779
rect 509 775 513 779
rect 517 775 521 779
rect 529 775 533 779
rect 537 775 541 779
rect 609 777 613 781
rect 633 777 637 781
rect 644 777 648 781
rect 654 777 658 781
rect 13 761 17 765
rect 400 769 404 773
rect 408 769 412 773
rect 580 769 584 773
rect 588 769 592 773
rect 14 725 18 729
rect 14 716 18 720
rect 14 708 18 712
rect 14 700 18 704
rect 14 688 18 692
rect 14 680 18 684
rect 124 657 128 661
rect 132 657 136 661
rect 144 657 148 661
rect 152 657 156 661
rect 304 657 308 661
rect 312 657 316 661
rect 324 657 328 661
rect 332 657 336 661
rect 657 659 661 663
rect 665 659 669 663
rect 677 659 681 663
rect 685 659 689 663
rect 837 659 841 663
rect 845 659 849 663
rect 857 659 861 663
rect 865 659 869 663
rect 14 641 18 645
rect 14 632 18 636
rect 62 634 66 638
rect 70 634 74 638
rect 82 634 86 638
rect 90 634 94 638
rect 182 647 186 651
rect 190 647 194 651
rect 202 647 206 651
rect 210 647 214 651
rect 14 624 18 628
rect 14 616 18 620
rect 14 604 18 608
rect 242 634 246 638
rect 250 634 254 638
rect 262 634 266 638
rect 270 634 274 638
rect 362 647 366 651
rect 370 647 374 651
rect 382 647 386 651
rect 390 647 394 651
rect 124 608 128 612
rect 132 608 136 612
rect 144 608 148 612
rect 595 636 599 640
rect 603 636 607 640
rect 615 636 619 640
rect 623 636 627 640
rect 715 649 719 653
rect 723 649 727 653
rect 735 649 739 653
rect 743 649 747 653
rect 152 608 156 612
rect 304 608 308 612
rect 312 608 316 612
rect 324 608 328 612
rect 775 636 779 640
rect 783 636 787 640
rect 795 636 799 640
rect 803 636 807 640
rect 895 649 899 653
rect 903 649 907 653
rect 915 649 919 653
rect 923 649 927 653
rect 332 608 336 612
rect 405 610 409 614
rect 429 610 433 614
rect 440 610 444 614
rect 450 610 454 614
rect 657 610 661 614
rect 665 610 669 614
rect 677 610 681 614
rect 685 610 689 614
rect 837 610 841 614
rect 845 610 849 614
rect 857 610 861 614
rect 865 610 869 614
rect 937 612 941 616
rect 961 612 965 616
rect 972 612 976 616
rect 982 612 986 616
rect 14 596 18 600
rect 195 602 199 606
rect 203 602 207 606
rect 375 602 379 606
rect 383 602 387 606
rect 728 604 732 608
rect 736 604 740 608
rect 908 604 912 608
rect 916 604 920 608
rect 14 554 18 558
rect 14 545 18 549
rect 14 537 18 541
rect 14 529 18 533
rect 14 517 18 521
rect 14 509 18 513
rect 315 502 319 506
rect 323 502 327 506
rect 335 502 339 506
rect 343 502 347 506
rect 495 502 499 506
rect 503 502 507 506
rect 515 502 519 506
rect 523 502 527 506
rect 253 479 257 483
rect 261 479 265 483
rect 273 479 277 483
rect 281 479 285 483
rect 373 492 377 496
rect 381 492 385 496
rect 393 492 397 496
rect 401 492 405 496
rect 15 466 19 470
rect 15 457 19 461
rect 433 479 437 483
rect 441 479 445 483
rect 453 479 457 483
rect 461 479 465 483
rect 553 492 557 496
rect 561 492 565 496
rect 573 492 577 496
rect 581 492 585 496
rect 315 453 319 457
rect 15 449 19 453
rect 323 453 327 457
rect 335 453 339 457
rect 343 453 347 457
rect 495 453 499 457
rect 503 453 507 457
rect 515 453 519 457
rect 523 453 527 457
rect 595 455 599 459
rect 619 455 623 459
rect 630 455 634 459
rect 640 455 644 459
rect 15 441 19 445
rect 15 429 19 433
rect 386 447 390 451
rect 394 447 398 451
rect 566 447 570 451
rect 574 447 578 451
rect 15 421 19 425
rect 145 401 149 405
rect 153 401 157 405
rect 165 401 169 405
rect 173 401 177 405
rect 16 385 20 389
rect 16 376 20 380
rect 83 378 87 382
rect 91 378 95 382
rect 103 378 107 382
rect 111 378 115 382
rect 203 391 207 395
rect 211 391 215 395
rect 223 391 227 395
rect 231 391 235 395
rect 16 368 20 372
rect 16 360 20 364
rect 16 348 20 352
rect 562 367 566 371
rect 570 367 574 371
rect 582 367 586 371
rect 590 367 594 371
rect 742 367 746 371
rect 750 367 754 371
rect 762 367 766 371
rect 770 367 774 371
rect 145 352 149 356
rect 153 352 157 356
rect 165 352 169 356
rect 173 352 177 356
rect 16 340 20 344
rect 216 346 220 350
rect 224 346 228 350
rect 500 344 504 348
rect 508 344 512 348
rect 520 344 524 348
rect 528 344 532 348
rect 620 357 624 361
rect 628 357 632 361
rect 640 357 644 361
rect 648 357 652 361
rect 680 344 684 348
rect 688 344 692 348
rect 700 344 704 348
rect 708 344 712 348
rect 800 357 804 361
rect 808 357 812 361
rect 820 357 824 361
rect 828 357 832 361
rect 562 318 566 322
rect 570 318 574 322
rect 582 318 586 322
rect 590 318 594 322
rect 742 318 746 322
rect 750 318 754 322
rect 762 318 766 322
rect 770 318 774 322
rect 842 320 846 324
rect 866 320 870 324
rect 877 320 881 324
rect 887 320 891 324
rect 16 301 20 305
rect 16 292 20 296
rect 633 312 637 316
rect 641 312 645 316
rect 813 312 817 316
rect 821 312 825 316
rect 16 284 20 288
rect 16 276 20 280
rect 16 264 20 268
rect 16 256 20 260
rect 16 214 20 218
rect 162 215 166 219
rect 170 215 174 219
rect 182 215 186 219
rect 190 215 194 219
rect 342 215 346 219
rect 350 215 354 219
rect 362 215 366 219
rect 370 215 374 219
rect 16 205 20 209
rect 16 197 20 201
rect 16 189 20 193
rect 16 177 20 181
rect 100 192 104 196
rect 108 192 112 196
rect 120 192 124 196
rect 128 192 132 196
rect 220 205 224 209
rect 228 205 232 209
rect 240 205 244 209
rect 248 205 252 209
rect 16 169 20 173
rect 280 192 284 196
rect 288 192 292 196
rect 300 192 304 196
rect 308 192 312 196
rect 400 205 404 209
rect 408 205 412 209
rect 420 205 424 209
rect 428 205 432 209
rect 162 166 166 170
rect 170 166 174 170
rect 182 166 186 170
rect 190 166 194 170
rect 342 166 346 170
rect 350 166 354 170
rect 362 166 366 170
rect 370 166 374 170
rect 442 168 446 172
rect 466 168 470 172
rect 477 168 481 172
rect 487 168 491 172
rect 585 168 589 172
rect 593 168 597 172
rect 605 168 609 172
rect 613 168 617 172
rect 765 168 769 172
rect 773 168 777 172
rect 785 168 789 172
rect 793 168 797 172
rect 233 160 237 164
rect 241 160 245 164
rect 413 160 417 164
rect 421 160 425 164
rect 523 145 527 149
rect 531 145 535 149
rect 543 145 547 149
rect 551 145 555 149
rect 643 158 647 162
rect 651 158 655 162
rect 663 158 667 162
rect 671 158 675 162
rect 17 126 21 130
rect 703 145 707 149
rect 711 145 715 149
rect 723 145 727 149
rect 731 145 735 149
rect 823 158 827 162
rect 831 158 835 162
rect 843 158 847 162
rect 851 158 855 162
rect 17 117 21 121
rect 585 119 589 123
rect 593 119 597 123
rect 605 119 609 123
rect 613 119 617 123
rect 765 119 769 123
rect 773 119 777 123
rect 785 119 789 123
rect 793 119 797 123
rect 865 121 869 125
rect 889 121 893 125
rect 900 121 904 125
rect 910 121 914 125
rect 17 109 21 113
rect 17 101 21 105
rect 17 89 21 93
rect 656 113 660 117
rect 664 113 668 117
rect 836 113 840 117
rect 844 113 848 117
rect 17 81 21 85
rect 18 45 22 49
rect 18 36 22 40
rect 18 28 22 32
rect 18 20 22 24
rect 18 8 22 12
rect 18 0 22 4
<< m2contact >>
rect 0 1259 4 1263
rect 26 1242 30 1246
rect 87 1259 91 1263
rect 131 1259 135 1263
rect 315 1260 319 1264
rect 359 1260 363 1264
rect 56 1243 60 1247
rect 87 1236 91 1240
rect 124 1220 128 1224
rect 131 1210 135 1214
rect 77 1193 81 1197
rect 115 1194 119 1198
rect 40 1172 44 1176
rect 27 1154 31 1158
rect 315 1237 319 1241
rect 352 1221 356 1225
rect 359 1211 363 1215
rect 305 1194 309 1198
rect 343 1195 347 1199
rect 203 1186 207 1190
rect 296 1188 301 1192
rect 431 1187 435 1191
rect 451 1185 456 1190
rect 77 1171 81 1175
rect 125 1171 129 1175
rect 305 1172 309 1176
rect 353 1172 357 1176
rect 70 1156 74 1160
rect 28 1073 32 1077
rect 2 1005 6 1009
rect 28 989 32 993
rect 74 1005 78 1009
rect 118 1005 122 1009
rect 254 1005 258 1009
rect 298 1005 302 1009
rect 58 989 62 993
rect 74 982 78 986
rect 214 974 218 978
rect 111 966 115 970
rect 118 956 122 960
rect 64 939 68 943
rect 102 940 106 944
rect 56 933 60 937
rect 238 989 242 993
rect 254 982 258 986
rect 394 976 398 980
rect 291 966 295 970
rect 235 946 240 951
rect 190 932 194 936
rect 298 956 302 960
rect 244 939 248 943
rect 282 940 286 944
rect 209 931 213 935
rect 569 1002 573 1006
rect 613 1002 617 1006
rect 560 986 565 991
rect 569 979 573 983
rect 606 963 610 967
rect 370 932 374 936
rect 397 931 401 935
rect 613 953 617 957
rect 559 936 563 940
rect 597 937 601 941
rect 29 902 33 906
rect 64 917 68 921
rect 112 917 116 921
rect 244 917 248 921
rect 292 917 296 921
rect 220 906 224 910
rect 397 906 401 910
rect 551 930 555 934
rect 685 929 689 933
rect 469 900 475 906
rect 559 914 563 918
rect 607 914 611 918
rect 3 833 8 838
rect 29 814 33 818
rect 277 834 281 838
rect 321 834 325 838
rect 457 834 461 838
rect 501 834 505 838
rect 277 811 281 815
rect 417 803 421 807
rect 314 795 318 799
rect 321 785 325 789
rect 267 768 271 772
rect 305 769 309 773
rect 259 762 263 766
rect 441 818 445 822
rect 457 811 461 815
rect 596 806 600 810
rect 494 795 498 799
rect 438 775 443 780
rect 393 761 397 765
rect 501 785 505 789
rect 447 768 451 772
rect 485 769 489 773
rect 412 760 416 764
rect 573 761 577 765
rect 600 760 604 764
rect 31 734 35 738
rect 267 746 271 750
rect 315 746 319 750
rect 447 746 451 750
rect 495 746 499 750
rect 423 735 427 739
rect 600 735 604 739
rect 816 691 820 695
rect 640 683 645 688
rect 5 666 9 670
rect 31 650 35 654
rect 72 667 76 671
rect 116 667 120 671
rect 252 667 256 671
rect 296 667 300 671
rect 55 651 59 655
rect 72 644 76 648
rect 212 636 216 640
rect 109 628 113 632
rect 116 618 120 622
rect 62 601 66 605
rect 100 602 104 606
rect 54 595 58 599
rect 235 651 239 655
rect 252 644 256 648
rect 392 636 396 640
rect 289 628 293 632
rect 233 608 238 613
rect 188 594 192 598
rect 296 618 300 622
rect 242 601 246 605
rect 280 602 284 606
rect 207 593 211 597
rect 605 669 609 673
rect 649 669 653 673
rect 785 669 789 673
rect 829 669 833 673
rect 639 653 643 657
rect 605 646 609 650
rect 745 638 749 642
rect 642 630 646 634
rect 368 594 372 598
rect 395 593 399 597
rect 649 620 653 624
rect 595 603 599 607
rect 633 604 637 608
rect 587 597 591 601
rect 43 579 47 583
rect 62 579 66 583
rect 110 579 114 583
rect 31 563 35 567
rect 242 579 246 583
rect 290 579 294 583
rect 218 568 222 572
rect 395 568 399 572
rect 816 654 820 658
rect 785 646 789 650
rect 822 630 826 634
rect 766 610 771 615
rect 721 596 725 600
rect 829 620 833 624
rect 775 603 779 607
rect 813 604 817 608
rect 740 595 744 599
rect 901 596 905 600
rect 928 595 932 599
rect 595 581 599 585
rect 643 581 647 585
rect 460 566 465 571
rect 775 581 779 585
rect 823 581 827 585
rect 751 570 755 574
rect 928 570 932 574
rect 263 512 267 516
rect 307 512 311 516
rect 443 512 447 516
rect 487 512 491 516
rect 31 474 35 478
rect 246 496 250 500
rect 263 489 267 493
rect 403 481 407 485
rect 300 473 304 477
rect 307 463 311 467
rect 253 446 257 450
rect 291 447 295 451
rect 245 439 249 443
rect 427 496 431 500
rect 443 489 447 493
rect 582 481 586 485
rect 480 473 484 477
rect 424 453 429 458
rect 379 439 383 443
rect 487 463 491 467
rect 433 446 437 450
rect 471 447 475 451
rect 398 438 402 442
rect 559 439 563 443
rect 586 438 590 442
rect 253 424 257 428
rect 301 424 305 428
rect 433 424 437 428
rect 481 424 485 428
rect 6 411 10 415
rect 32 394 36 398
rect 93 411 97 415
rect 137 411 141 415
rect 409 413 413 417
rect 586 413 590 417
rect 58 394 62 398
rect 93 388 97 392
rect 232 382 236 386
rect 130 372 134 376
rect 137 362 141 366
rect 83 345 87 349
rect 121 346 125 350
rect 640 402 644 406
rect 722 390 726 394
rect 510 377 514 381
rect 554 377 558 381
rect 690 377 694 381
rect 734 377 738 381
rect 46 323 50 327
rect 32 309 36 313
rect 541 361 545 365
rect 209 338 213 342
rect 273 336 278 342
rect 510 354 514 358
rect 650 346 654 350
rect 547 338 551 342
rect 83 323 87 327
rect 131 323 135 327
rect 76 310 80 314
rect 472 305 478 311
rect 554 328 558 332
rect 500 311 504 315
rect 538 312 542 316
rect 721 361 725 365
rect 690 354 694 358
rect 727 338 731 342
rect 671 318 676 323
rect 626 304 630 308
rect 734 328 738 332
rect 680 311 684 315
rect 718 312 722 316
rect 645 303 649 307
rect 806 304 810 308
rect 833 303 837 307
rect 500 289 504 293
rect 548 289 552 293
rect 680 289 684 293
rect 728 289 732 293
rect 656 278 660 282
rect 833 278 837 282
rect 697 256 702 261
rect 6 234 10 238
rect 32 223 36 227
rect 73 224 77 228
rect 110 225 114 229
rect 154 225 158 229
rect 290 225 294 229
rect 334 225 338 229
rect 110 202 114 206
rect 250 194 254 198
rect 147 186 151 190
rect 33 135 37 139
rect 154 176 158 180
rect 100 159 104 163
rect 138 160 142 164
rect 273 209 277 213
rect 290 202 294 206
rect 429 197 433 201
rect 327 186 331 190
rect 271 166 276 171
rect 226 152 230 156
rect 334 176 338 180
rect 280 159 284 163
rect 318 160 322 164
rect 245 151 249 155
rect 533 178 537 182
rect 577 178 581 182
rect 713 178 717 182
rect 757 178 761 182
rect 406 152 410 156
rect 433 151 437 155
rect 533 155 537 159
rect 673 147 677 151
rect 73 136 77 140
rect 100 137 104 141
rect 148 137 152 141
rect 280 137 284 141
rect 328 137 332 141
rect 570 139 574 143
rect 256 126 260 130
rect 433 126 437 130
rect 577 129 581 133
rect 523 112 527 116
rect 561 113 565 117
rect 515 106 519 110
rect 697 162 701 166
rect 713 155 717 159
rect 750 139 754 143
rect 694 119 699 124
rect 649 105 653 109
rect 757 129 761 133
rect 703 112 707 116
rect 741 113 745 117
rect 668 104 672 108
rect 829 105 833 109
rect 856 104 860 108
rect 523 90 527 94
rect 571 90 575 94
rect 703 90 707 94
rect 751 90 755 94
rect 33 54 37 58
rect 679 79 683 83
rect 856 79 860 83
<< psubstratepcontact >>
rect 39 1311 43 1315
rect 39 1276 43 1280
rect 39 1224 43 1228
rect 139 1220 143 1224
rect 367 1221 371 1225
rect 39 1189 43 1193
rect 99 1171 103 1175
rect 139 1171 143 1175
rect 167 1171 171 1175
rect 196 1171 200 1175
rect 219 1170 223 1174
rect 327 1172 331 1176
rect 367 1172 371 1176
rect 395 1172 399 1176
rect 424 1172 428 1176
rect 447 1171 451 1175
rect 40 1136 44 1140
rect 40 1101 44 1105
rect 41 1055 45 1059
rect 41 1020 45 1024
rect 41 971 45 975
rect 126 966 130 970
rect 306 966 310 970
rect 621 963 625 967
rect 41 936 45 940
rect 86 917 90 921
rect 126 917 130 921
rect 154 917 158 921
rect 183 917 187 921
rect 206 916 210 920
rect 266 917 270 921
rect 306 917 310 921
rect 334 917 338 921
rect 363 917 367 921
rect 386 916 390 920
rect 419 916 423 920
rect 581 914 585 918
rect 621 914 625 918
rect 649 914 653 918
rect 678 914 682 918
rect 701 913 705 917
rect 41 884 45 888
rect 41 849 45 853
rect 42 796 46 800
rect 329 795 333 799
rect 509 795 513 799
rect 42 761 46 765
rect 289 746 293 750
rect 329 746 333 750
rect 357 746 361 750
rect 386 746 390 750
rect 409 745 413 749
rect 469 746 473 750
rect 509 746 513 750
rect 537 746 541 750
rect 566 746 570 750
rect 589 745 593 749
rect 621 745 625 749
rect 43 715 47 719
rect 43 680 47 684
rect 43 631 47 635
rect 124 628 128 632
rect 304 628 308 632
rect 657 630 661 634
rect 837 630 841 634
rect 43 596 47 600
rect 84 579 88 583
rect 124 579 128 583
rect 152 579 156 583
rect 181 579 185 583
rect 204 578 208 582
rect 264 579 268 583
rect 304 579 308 583
rect 332 579 336 583
rect 361 579 365 583
rect 384 578 388 582
rect 417 578 421 582
rect 617 581 621 585
rect 657 581 661 585
rect 685 581 689 585
rect 714 581 718 585
rect 737 580 741 584
rect 797 581 801 585
rect 837 581 841 585
rect 865 581 869 585
rect 894 581 898 585
rect 917 580 921 584
rect 949 580 953 584
rect 43 544 47 548
rect 43 509 47 513
rect 44 456 48 460
rect 315 473 319 477
rect 495 473 499 477
rect 44 421 48 425
rect 275 424 279 428
rect 315 424 319 428
rect 343 424 347 428
rect 372 424 376 428
rect 395 423 399 427
rect 455 424 459 428
rect 495 424 499 428
rect 523 424 527 428
rect 552 424 556 428
rect 575 423 579 427
rect 607 423 611 427
rect 45 375 49 379
rect 145 372 149 376
rect 45 340 49 344
rect 105 323 109 327
rect 145 323 149 327
rect 173 323 177 327
rect 202 323 206 327
rect 225 322 229 326
rect 562 338 566 342
rect 742 338 746 342
rect 45 291 49 295
rect 522 289 526 293
rect 562 289 566 293
rect 590 289 594 293
rect 619 289 623 293
rect 642 288 646 292
rect 702 289 706 293
rect 742 289 746 293
rect 770 289 774 293
rect 799 289 803 293
rect 822 288 826 292
rect 854 288 858 292
rect 45 256 49 260
rect 45 204 49 208
rect 45 169 49 173
rect 162 186 166 190
rect 342 186 346 190
rect 122 137 126 141
rect 162 137 166 141
rect 190 137 194 141
rect 219 137 223 141
rect 242 136 246 140
rect 302 137 306 141
rect 342 137 346 141
rect 370 137 374 141
rect 399 137 403 141
rect 422 136 426 140
rect 454 136 458 140
rect 585 139 589 143
rect 46 116 50 120
rect 765 139 769 143
rect 545 90 549 94
rect 585 90 589 94
rect 613 90 617 94
rect 642 90 646 94
rect 665 89 669 93
rect 725 90 729 94
rect 765 90 769 94
rect 793 90 797 94
rect 822 90 826 94
rect 845 89 849 93
rect 877 89 881 93
rect 46 81 50 85
rect 47 35 51 39
rect 47 0 51 4
<< nsubstratencontact >>
rect 0 1312 4 1316
rect 0 1296 4 1300
rect 0 1276 4 1280
rect 139 1259 143 1263
rect 159 1259 163 1263
rect 197 1259 201 1263
rect 367 1260 371 1264
rect 387 1260 391 1264
rect 425 1260 429 1264
rect 197 1249 201 1253
rect 217 1249 221 1253
rect 425 1250 429 1254
rect 445 1250 449 1254
rect 77 1236 81 1240
rect 97 1236 101 1240
rect 0 1225 4 1229
rect 0 1209 4 1213
rect 305 1237 309 1241
rect 325 1237 329 1241
rect 139 1210 143 1214
rect 159 1210 163 1214
rect 221 1204 225 1208
rect 367 1211 371 1215
rect 387 1211 391 1215
rect 449 1205 453 1209
rect 0 1189 4 1193
rect 1 1137 5 1141
rect 1 1121 5 1125
rect 1 1101 5 1105
rect 2 1056 6 1060
rect 2 1040 6 1044
rect 2 1020 6 1024
rect 126 1005 130 1009
rect 146 1005 150 1009
rect 184 1005 188 1009
rect 306 1005 310 1009
rect 326 1005 330 1009
rect 364 1005 368 1009
rect 621 1002 625 1006
rect 641 1002 645 1006
rect 679 1002 683 1006
rect 184 995 188 999
rect 204 995 208 999
rect 364 995 368 999
rect 384 995 388 999
rect 64 982 68 986
rect 84 982 88 986
rect 2 972 6 976
rect 2 956 6 960
rect 244 982 248 986
rect 264 982 268 986
rect 679 992 683 996
rect 699 992 703 996
rect 126 956 130 960
rect 146 956 150 960
rect 208 950 212 954
rect 559 979 563 983
rect 579 979 583 983
rect 306 956 310 960
rect 326 956 330 960
rect 407 957 411 961
rect 442 957 446 961
rect 388 950 392 954
rect 621 953 625 957
rect 641 953 645 957
rect 2 936 6 940
rect 703 947 707 951
rect 2 885 6 889
rect 2 869 6 873
rect 2 849 6 853
rect 329 834 333 838
rect 349 834 353 838
rect 387 834 391 838
rect 509 834 513 838
rect 529 834 533 838
rect 567 834 571 838
rect 387 824 391 828
rect 407 824 411 828
rect 567 824 571 828
rect 587 824 591 828
rect 267 811 271 815
rect 287 811 291 815
rect 3 797 7 801
rect 3 781 7 785
rect 447 811 451 815
rect 467 811 471 815
rect 329 785 333 789
rect 349 785 353 789
rect 411 779 415 783
rect 509 785 513 789
rect 529 785 533 789
rect 609 786 613 790
rect 644 786 648 790
rect 591 779 595 783
rect 3 761 7 765
rect 4 716 8 720
rect 4 700 8 704
rect 4 680 8 684
rect 124 667 128 671
rect 144 667 148 671
rect 182 667 186 671
rect 304 667 308 671
rect 324 667 328 671
rect 362 667 366 671
rect 657 669 661 673
rect 677 669 681 673
rect 715 669 719 673
rect 837 669 841 673
rect 857 669 861 673
rect 895 669 899 673
rect 182 657 186 661
rect 202 657 206 661
rect 362 657 366 661
rect 382 657 386 661
rect 715 659 719 663
rect 735 659 739 663
rect 895 659 899 663
rect 915 659 919 663
rect 62 644 66 648
rect 82 644 86 648
rect 4 632 8 636
rect 4 616 8 620
rect 242 644 246 648
rect 262 644 266 648
rect 595 646 599 650
rect 615 646 619 650
rect 124 618 128 622
rect 144 618 148 622
rect 206 612 210 616
rect 304 618 308 622
rect 324 618 328 622
rect 405 619 409 623
rect 440 619 444 623
rect 386 612 390 616
rect 775 646 779 650
rect 795 646 799 650
rect 657 620 661 624
rect 677 620 681 624
rect 739 614 743 618
rect 837 620 841 624
rect 857 620 861 624
rect 937 621 941 625
rect 972 621 976 625
rect 919 614 923 618
rect 4 596 8 600
rect 4 545 8 549
rect 4 529 8 533
rect 4 509 8 513
rect 315 512 319 516
rect 335 512 339 516
rect 373 512 377 516
rect 495 512 499 516
rect 515 512 519 516
rect 553 512 557 516
rect 373 502 377 506
rect 393 502 397 506
rect 553 502 557 506
rect 573 502 577 506
rect 253 489 257 493
rect 273 489 277 493
rect 5 457 9 461
rect 433 489 437 493
rect 453 489 457 493
rect 315 463 319 467
rect 335 463 339 467
rect 397 457 401 461
rect 495 463 499 467
rect 515 463 519 467
rect 595 464 599 468
rect 630 464 634 468
rect 577 457 581 461
rect 5 441 9 445
rect 5 421 9 425
rect 145 411 149 415
rect 165 411 169 415
rect 203 411 207 415
rect 203 401 207 405
rect 223 401 227 405
rect 83 388 87 392
rect 103 388 107 392
rect 6 376 10 380
rect 6 360 10 364
rect 562 377 566 381
rect 582 377 586 381
rect 620 377 624 381
rect 742 377 746 381
rect 762 377 766 381
rect 800 377 804 381
rect 620 367 624 371
rect 640 367 644 371
rect 800 367 804 371
rect 820 367 824 371
rect 145 362 149 366
rect 165 362 169 366
rect 227 356 231 360
rect 500 354 504 358
rect 520 354 524 358
rect 6 340 10 344
rect 680 354 684 358
rect 700 354 704 358
rect 562 328 566 332
rect 582 328 586 332
rect 644 322 648 326
rect 742 328 746 332
rect 762 328 766 332
rect 842 329 846 333
rect 877 329 881 333
rect 824 322 828 326
rect 6 292 10 296
rect 6 276 10 280
rect 6 256 10 260
rect 162 225 166 229
rect 182 225 186 229
rect 220 225 224 229
rect 342 225 346 229
rect 362 225 366 229
rect 400 225 404 229
rect 220 215 224 219
rect 240 215 244 219
rect 400 215 404 219
rect 420 215 424 219
rect 6 205 10 209
rect 100 202 104 206
rect 120 202 124 206
rect 6 189 10 193
rect 6 169 10 173
rect 280 202 284 206
rect 300 202 304 206
rect 162 176 166 180
rect 182 176 186 180
rect 244 170 248 174
rect 342 176 346 180
rect 362 176 366 180
rect 442 177 446 181
rect 477 177 481 181
rect 585 178 589 182
rect 605 178 609 182
rect 643 178 647 182
rect 765 178 769 182
rect 785 178 789 182
rect 823 178 827 182
rect 424 170 428 174
rect 643 168 647 172
rect 663 168 667 172
rect 823 168 827 172
rect 843 168 847 172
rect 523 155 527 159
rect 543 155 547 159
rect 703 155 707 159
rect 723 155 727 159
rect 585 129 589 133
rect 605 129 609 133
rect 7 117 11 121
rect 667 123 671 127
rect 765 129 769 133
rect 785 129 789 133
rect 865 130 869 134
rect 900 130 904 134
rect 847 123 851 127
rect 7 101 11 105
rect 7 81 11 85
rect 8 36 12 40
rect 8 20 12 24
rect 8 0 12 4
<< labels >>
rlabel metal1 11 11 11 11 7 Vdd
rlabel metal1 50 11 50 11 7 Gnd
rlabel metal1 10 92 10 92 7 Vdd
rlabel metal1 49 92 49 92 7 Gnd
rlabel metal1 9 180 9 180 7 Vdd
rlabel metal1 48 180 48 180 7 Gnd
rlabel metal1 9 267 9 267 7 Vdd
rlabel metal1 48 267 48 267 7 Gnd
rlabel metal1 9 351 9 351 7 Vdd
rlabel metal1 48 351 48 351 7 Gnd
rlabel metal1 8 432 8 432 7 Vdd
rlabel metal1 47 432 47 432 7 Gnd
rlabel metal1 7 520 7 520 7 Vdd
rlabel metal1 46 520 46 520 7 Gnd
rlabel metal1 7 607 7 607 7 Vdd
rlabel metal1 46 607 46 607 7 Gnd
rlabel metal1 7 691 7 691 7 Vdd
rlabel metal1 46 691 46 691 7 Gnd
rlabel metal1 6 772 6 772 7 Vdd
rlabel metal1 45 772 45 772 7 Gnd
rlabel metal1 5 860 5 860 7 Vdd
rlabel metal1 44 860 44 860 7 Gnd
rlabel metal1 5 947 5 947 7 Vdd
rlabel metal1 44 947 44 947 7 Gnd
rlabel metal1 5 1031 5 1031 7 Vdd
rlabel metal1 44 1031 44 1031 7 Gnd
rlabel metal1 4 1112 4 1112 7 Vdd
rlabel metal1 43 1112 43 1112 7 Gnd
rlabel metal1 3 1200 3 1200 7 Vdd
rlabel metal1 42 1200 42 1200 7 Gnd
rlabel metal1 3 1287 3 1287 7 Vdd
rlabel metal1 42 1287 42 1287 7 Gnd
rlabel metal1 32 46 32 46 7 x3y3
rlabel metal1 30 302 30 302 1 x2y2
rlabel metal1 30 386 30 386 1 x1y3
rlabel metal1 29 467 29 467 1 x3y1
rlabel metal1 26 1066 26 1066 1 x2y0
rlabel metal1 25 1147 25 1147 1 x1y0
rlabel metal1 24 1235 24 1235 1 x0y1
rlabel metal1 115 325 115 325 1 Gnd
rlabel metal1 118 412 118 412 1 Vdd
rlabel metal1 78 396 78 396 3 P13
rlabel metal1 78 340 78 340 3 P22
rlabel metal1 31 127 31 127 1 x2y3
rlabel metal1 30 215 30 215 1 x3y2
rlabel metal1 28 555 28 555 1 x2y1
rlabel metal1 28 642 28 642 1 x1y2
rlabel metal1 28 726 28 726 1 x0y3
rlabel metal1 27 807 27 807 1 x3y0
rlabel metal1 26 895 26 895 1 x0y2
rlabel metal1 26 982 26 982 1 x1y1
rlabel metal1 228 339 228 339 3 C04
rlabel metal1 312 139 312 139 1 Gnd
rlabel metal1 315 226 315 226 1 Vdd
rlabel metal1 132 139 132 139 1 Gnd
rlabel metal1 135 226 135 226 1 Vdd
rlabel metal1 449 139 449 139 3 Gnd
rlabel metal1 460 179 460 179 1 Vdd
rlabel metal1 95 210 95 210 3 P23
rlabel polycontact 104 187 104 187 3 P23
rlabel metal1 95 154 95 154 3 P32
rlabel polycontact 124 180 124 180 3 P32
rlabel polycontact 166 210 166 210 3 P23
rlabel polycontact 186 154 186 154 3 P32
rlabel metal1 109 1173 109 1173 1 Gnd
rlabel metal1 112 1260 112 1260 1 Vdd
rlabel metal1 72 1244 72 1244 3 P01
rlabel metal1 72 1188 72 1188 3 P10
rlabel metal1 222 1187 222 1187 3 C01
rlabel metal1 227 1234 227 1234 1 S01
rlabel metal1 276 919 276 919 1 Gnd
rlabel metal1 279 1006 279 1006 1 Vdd
rlabel metal1 96 919 96 919 1 Gnd
rlabel metal1 99 1006 99 1006 1 Vdd
rlabel metal1 59 987 59 987 5 P11
rlabel metal1 59 939 59 939 1 P02
rlabel polycontact 68 967 68 967 1 P11
rlabel polycontact 130 990 130 990 1 P11
rlabel polycontact 88 960 88 960 1 P02
rlabel polycontact 150 934 150 934 1 P02
rlabel metal1 239 987 239 987 3 P20
rlabel metal1 274 581 274 581 1 Gnd
rlabel metal1 277 668 277 668 1 Vdd
rlabel metal1 94 581 94 581 1 Gnd
rlabel metal1 97 668 97 668 1 Vdd
rlabel metal1 57 648 57 648 1 P12
rlabel metal1 57 601 57 601 1 P21
rlabel polycontact 148 596 148 596 1 P21
rlabel polycontact 86 622 86 622 1 P21
rlabel polycontact 66 629 66 629 1 P12
rlabel polycontact 128 652 128 652 1 P12
rlabel metal1 237 649 237 649 1 P03
rlabel metal1 337 1174 337 1174 1 Gnd
rlabel metal1 340 1261 340 1261 1 Vdd
rlabel metal1 300 1245 300 1245 1 C01
rlabel polycontact 309 1222 309 1222 1 C01
rlabel polycontact 371 1245 371 1245 1 C01
rlabel metal1 455 1235 455 1235 1 S11
rlabel polycontact 391 1189 391 1189 1 S02
rlabel polycontact 329 1215 329 1215 1 S02
rlabel metal1 414 919 414 919 3 Gnd
rlabel metal1 425 959 425 959 1 Vdd
rlabel metal1 455 937 455 937 1 C02
rlabel metal1 393 980 393 980 1 S02
rlabel metal1 300 1193 300 1193 1 S02
rlabel metal1 479 748 479 748 1 Gnd
rlabel metal1 482 835 482 835 1 Vdd
rlabel metal1 299 748 299 748 1 Gnd
rlabel metal1 302 835 302 835 1 Vdd
rlabel metal1 616 748 616 748 3 Gnd
rlabel metal1 627 788 627 788 1 Vdd
rlabel polycontact 333 819 333 819 1 in_1
rlabel polycontact 353 763 353 763 1 in_2
rlabel polycontact 291 789 291 789 1 in_2
rlabel polycontact 271 796 271 796 1 in_1
rlabel metal1 262 820 262 820 3 P30
rlabel metal1 262 767 262 767 1 S03
rlabel metal1 412 581 412 581 3 Gnd
rlabel metal1 423 621 423 621 1 Vdd
rlabel metal1 392 642 392 642 1 S03
rlabel metal1 453 599 453 599 1 C03
rlabel metal1 442 816 442 816 5 C02
rlabel metal1 657 766 657 766 1 C12
rlabel metal1 613 466 613 466 1 Vdd
rlabel metal1 602 426 602 426 3 Gnd
rlabel metal1 288 513 288 513 1 Vdd
rlabel metal1 285 426 285 426 1 Gnd
rlabel metal1 468 513 468 513 1 Vdd
rlabel metal1 465 426 465 426 1 Gnd
rlabel metal1 253 497 253 497 1 P31
rlabel polycontact 257 474 257 474 1 P31
rlabel polycontact 319 497 319 497 1 P31
rlabel metal1 429 493 429 493 1 C03
rlabel metal1 583 487 583 487 1 S13
rlabel metal1 643 444 643 444 1 C13
rlabel metal1 248 444 248 444 1 S04
rlabel polycontact 339 441 339 441 1 S04
rlabel polycontact 277 467 277 467 1 S04
rlabel metal1 231 386 231 386 7 S04
rlabel metal1 735 92 735 92 1 Gnd
rlabel metal1 738 179 738 179 1 Vdd
rlabel metal1 555 92 555 92 1 Gnd
rlabel metal1 558 179 558 179 1 Vdd
rlabel metal1 872 92 872 92 3 Gnd
rlabel metal1 913 110 913 110 1 C_out
rlabel metal1 883 132 883 132 1 Vdd
rlabel metal1 490 157 490 157 1 C14
rlabel metal1 518 163 518 163 1 C14
rlabel polycontact 589 163 589 163 1 C14
rlabel polycontact 527 140 527 140 1 C14
rlabel metal1 698 158 698 158 1 C23
rlabel metal1 853 153 853 153 1 S24
rlabel metal1 518 112 518 112 1 P33
rlabel polycontact 547 133 547 133 1 P33
rlabel polycontact 609 107 609 107 1 P33
rlabel metal1 712 291 712 291 1 Gnd
rlabel metal1 715 378 715 378 1 Vdd
rlabel metal1 532 291 532 291 1 Gnd
rlabel metal1 535 378 535 378 1 Vdd
rlabel metal1 849 291 849 291 3 Gnd
rlabel metal1 860 331 860 331 1 Vdd
rlabel metal1 890 309 890 309 1 C23
rlabel metal1 428 200 428 200 1 S14
rlabel metal1 495 306 495 306 1 S14
rlabel polycontact 586 306 586 306 1 S14
rlabel polycontact 524 332 524 332 1 S14
rlabel metal1 495 362 495 362 1 C13
rlabel polycontact 504 339 504 339 1 C13
rlabel polycontact 566 362 566 362 1 C13
rlabel metal1 830 352 830 352 1 S23
rlabel metal1 675 362 675 362 1 C22
rlabel metal1 593 809 593 809 1 S12
rlabel metal1 591 916 591 916 1 Gnd
rlabel metal1 594 1003 594 1003 1 Vdd
rlabel metal1 553 936 553 936 1 S12
rlabel polycontact 583 957 583 957 1 S12
rlabel polycontact 645 931 645 931 1 S12
rlabel metal1 704 930 704 930 1 C21
rlabel metal1 709 977 709 977 1 S21
rlabel polycontact 563 964 563 964 1 C11
rlabel polycontact 625 987 625 987 1 C11
rlabel metal1 554 985 554 985 1 C11
rlabel metal1 450 1190 450 1190 1 C11
rlabel metal1 807 583 807 583 1 Gnd
rlabel metal1 810 670 810 670 1 Vdd
rlabel metal1 627 583 627 583 1 Gnd
rlabel metal1 630 670 630 670 1 Vdd
rlabel metal1 944 583 944 583 3 Gnd
rlabel metal1 955 623 955 623 1 Vdd
rlabel metal1 590 602 590 602 1 S13
rlabel polycontact 681 598 681 598 1 S13
rlabel polycontact 619 624 619 624 1 S13
rlabel metal1 590 654 590 654 1 C12
rlabel polycontact 599 631 599 631 1 C12
rlabel polycontact 661 654 661 654 1 C12
rlabel metal1 925 644 925 644 1 S22
rlabel metal1 985 603 985 603 1 C22
rlabel metal1 770 654 770 654 1 C21
rlabel metal1 24 1322 24 1322 7 P00
rlabel polycontact 26 1300 26 1300 1 y0a
rlabel polycontact 19 1280 19 1280 1 x0a
rlabel polycontact 26 1213 26 1213 1 y1a
rlabel polycontact 19 1193 19 1193 1 x0b
rlabel polycontact 27 1125 27 1125 1 y0b
rlabel polycontact 20 1105 20 1105 1 x1a
rlabel polycontact 28 1044 28 1044 1 y0c
rlabel polycontact 21 1024 21 1024 1 x2a
rlabel polycontact 28 960 28 960 1 y1b
rlabel polycontact 21 940 21 940 1 x1b
rlabel polycontact 28 873 28 873 1 y2a
rlabel polycontact 21 853 21 853 1 x0c
rlabel polycontact 29 785 29 785 1 y0d
rlabel polycontact 22 765 22 765 1 x3a
rlabel polycontact 30 704 30 704 1 y3a
rlabel polycontact 23 684 23 684 1 x0d
rlabel polycontact 30 620 30 620 1 y2b
rlabel polycontact 23 600 23 600 1 x1c
rlabel polycontact 30 533 30 533 1 y1c
rlabel polycontact 23 513 23 513 1 x2b
rlabel polycontact 31 445 31 445 1 y1d
rlabel polycontact 24 425 24 425 1 x3b
rlabel polycontact 32 364 32 364 1 y3b
rlabel polycontact 25 344 25 344 1 x1d
rlabel polycontact 32 280 32 280 1 y2c
rlabel polycontact 25 260 25 260 1 x2c
rlabel polycontact 32 193 32 193 1 y2d
rlabel polycontact 25 173 25 173 1 x3c
rlabel polycontact 33 105 33 105 1 y3c
rlabel polycontact 26 85 26 85 1 x2d
rlabel polycontact 34 24 34 24 1 y3d
rlabel polycontact 27 4 27 4 1 x3d
<< end >>
